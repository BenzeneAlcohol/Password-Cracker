magic
tech sky130A
magscale 1 2
timestamp 1679563233
<< obsli1 >>
rect 1104 2159 85192 85969
<< obsm1 >>
rect 14 1572 86098 87440
<< metal2 >>
rect 662 87640 718 88440
rect 1950 87640 2006 88440
rect 3238 87640 3294 88440
rect 3882 87640 3938 88440
rect 5170 87640 5226 88440
rect 6458 87640 6514 88440
rect 7746 87640 7802 88440
rect 9034 87640 9090 88440
rect 9678 87640 9734 88440
rect 10966 87640 11022 88440
rect 12254 87640 12310 88440
rect 13542 87640 13598 88440
rect 14830 87640 14886 88440
rect 15474 87640 15530 88440
rect 16762 87640 16818 88440
rect 18050 87640 18106 88440
rect 19338 87640 19394 88440
rect 20626 87640 20682 88440
rect 21270 87640 21326 88440
rect 22558 87640 22614 88440
rect 23846 87640 23902 88440
rect 25134 87640 25190 88440
rect 26422 87640 26478 88440
rect 27066 87640 27122 88440
rect 28354 87640 28410 88440
rect 29642 87640 29698 88440
rect 30930 87640 30986 88440
rect 32218 87640 32274 88440
rect 33506 87640 33562 88440
rect 34150 87640 34206 88440
rect 35438 87640 35494 88440
rect 36726 87640 36782 88440
rect 38014 87640 38070 88440
rect 39302 87640 39358 88440
rect 39946 87640 40002 88440
rect 41234 87640 41290 88440
rect 42522 87640 42578 88440
rect 43810 87640 43866 88440
rect 45098 87640 45154 88440
rect 45742 87640 45798 88440
rect 47030 87640 47086 88440
rect 48318 87640 48374 88440
rect 49606 87640 49662 88440
rect 50894 87640 50950 88440
rect 51538 87640 51594 88440
rect 52826 87640 52882 88440
rect 54114 87640 54170 88440
rect 55402 87640 55458 88440
rect 56690 87640 56746 88440
rect 57334 87640 57390 88440
rect 58622 87640 58678 88440
rect 59910 87640 59966 88440
rect 61198 87640 61254 88440
rect 62486 87640 62542 88440
rect 63130 87640 63186 88440
rect 64418 87640 64474 88440
rect 65706 87640 65762 88440
rect 66994 87640 67050 88440
rect 68282 87640 68338 88440
rect 68926 87640 68982 88440
rect 70214 87640 70270 88440
rect 71502 87640 71558 88440
rect 72790 87640 72846 88440
rect 74078 87640 74134 88440
rect 74722 87640 74778 88440
rect 76010 87640 76066 88440
rect 77298 87640 77354 88440
rect 78586 87640 78642 88440
rect 79874 87640 79930 88440
rect 80518 87640 80574 88440
rect 81806 87640 81862 88440
rect 83094 87640 83150 88440
rect 84382 87640 84438 88440
rect 85670 87640 85726 88440
rect 18 0 74 800
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 38014 0 38070 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 49606 0 49662 800
rect 50894 0 50950 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 55402 0 55458 800
rect 56690 0 56746 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59910 0 59966 800
rect 61198 0 61254 800
rect 62486 0 62542 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66994 0 67050 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 77298 0 77354 800
rect 78586 0 78642 800
rect 79874 0 79930 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85670 0 85726 800
<< obsm2 >>
rect 20 87584 606 87825
rect 774 87584 1894 87825
rect 2062 87584 3182 87825
rect 3350 87584 3826 87825
rect 3994 87584 5114 87825
rect 5282 87584 6402 87825
rect 6570 87584 7690 87825
rect 7858 87584 8978 87825
rect 9146 87584 9622 87825
rect 9790 87584 10910 87825
rect 11078 87584 12198 87825
rect 12366 87584 13486 87825
rect 13654 87584 14774 87825
rect 14942 87584 15418 87825
rect 15586 87584 16706 87825
rect 16874 87584 17994 87825
rect 18162 87584 19282 87825
rect 19450 87584 20570 87825
rect 20738 87584 21214 87825
rect 21382 87584 22502 87825
rect 22670 87584 23790 87825
rect 23958 87584 25078 87825
rect 25246 87584 26366 87825
rect 26534 87584 27010 87825
rect 27178 87584 28298 87825
rect 28466 87584 29586 87825
rect 29754 87584 30874 87825
rect 31042 87584 32162 87825
rect 32330 87584 33450 87825
rect 33618 87584 34094 87825
rect 34262 87584 35382 87825
rect 35550 87584 36670 87825
rect 36838 87584 37958 87825
rect 38126 87584 39246 87825
rect 39414 87584 39890 87825
rect 40058 87584 41178 87825
rect 41346 87584 42466 87825
rect 42634 87584 43754 87825
rect 43922 87584 45042 87825
rect 45210 87584 45686 87825
rect 45854 87584 46974 87825
rect 47142 87584 48262 87825
rect 48430 87584 49550 87825
rect 49718 87584 50838 87825
rect 51006 87584 51482 87825
rect 51650 87584 52770 87825
rect 52938 87584 54058 87825
rect 54226 87584 55346 87825
rect 55514 87584 56634 87825
rect 56802 87584 57278 87825
rect 57446 87584 58566 87825
rect 58734 87584 59854 87825
rect 60022 87584 61142 87825
rect 61310 87584 62430 87825
rect 62598 87584 63074 87825
rect 63242 87584 64362 87825
rect 64530 87584 65650 87825
rect 65818 87584 66938 87825
rect 67106 87584 68226 87825
rect 68394 87584 68870 87825
rect 69038 87584 70158 87825
rect 70326 87584 71446 87825
rect 71614 87584 72734 87825
rect 72902 87584 74022 87825
rect 74190 87584 74666 87825
rect 74834 87584 75954 87825
rect 76122 87584 77242 87825
rect 77410 87584 78530 87825
rect 78698 87584 79818 87825
rect 79986 87584 80462 87825
rect 80630 87584 81750 87825
rect 81918 87584 83038 87825
rect 83206 87584 84326 87825
rect 84494 87584 85614 87825
rect 85782 87584 86092 87825
rect 20 856 86092 87584
rect 130 711 606 856
rect 774 711 1894 856
rect 2062 711 3182 856
rect 3350 711 4470 856
rect 4638 711 5758 856
rect 5926 711 6402 856
rect 6570 711 7690 856
rect 7858 711 8978 856
rect 9146 711 10266 856
rect 10434 711 11554 856
rect 11722 711 12198 856
rect 12366 711 13486 856
rect 13654 711 14774 856
rect 14942 711 16062 856
rect 16230 711 17350 856
rect 17518 711 17994 856
rect 18162 711 19282 856
rect 19450 711 20570 856
rect 20738 711 21858 856
rect 22026 711 23146 856
rect 23314 711 23790 856
rect 23958 711 25078 856
rect 25246 711 26366 856
rect 26534 711 27654 856
rect 27822 711 28942 856
rect 29110 711 29586 856
rect 29754 711 30874 856
rect 31042 711 32162 856
rect 32330 711 33450 856
rect 33618 711 34738 856
rect 34906 711 35382 856
rect 35550 711 36670 856
rect 36838 711 37958 856
rect 38126 711 39246 856
rect 39414 711 40534 856
rect 40702 711 41178 856
rect 41346 711 42466 856
rect 42634 711 43754 856
rect 43922 711 45042 856
rect 45210 711 46330 856
rect 46498 711 46974 856
rect 47142 711 48262 856
rect 48430 711 49550 856
rect 49718 711 50838 856
rect 51006 711 52126 856
rect 52294 711 52770 856
rect 52938 711 54058 856
rect 54226 711 55346 856
rect 55514 711 56634 856
rect 56802 711 57922 856
rect 58090 711 58566 856
rect 58734 711 59854 856
rect 60022 711 61142 856
rect 61310 711 62430 856
rect 62598 711 63718 856
rect 63886 711 64362 856
rect 64530 711 65650 856
rect 65818 711 66938 856
rect 67106 711 68226 856
rect 68394 711 69514 856
rect 69682 711 70158 856
rect 70326 711 71446 856
rect 71614 711 72734 856
rect 72902 711 74022 856
rect 74190 711 75310 856
rect 75478 711 75954 856
rect 76122 711 77242 856
rect 77410 711 78530 856
rect 78698 711 79818 856
rect 79986 711 81106 856
rect 81274 711 81750 856
rect 81918 711 83038 856
rect 83206 711 84326 856
rect 84494 711 85614 856
rect 85782 711 86092 856
<< metal3 >>
rect 0 87728 800 87848
rect 85496 87728 86296 87848
rect 0 86368 800 86488
rect 85496 86368 86296 86488
rect 0 85688 800 85808
rect 85496 85008 86296 85128
rect 0 84328 800 84448
rect 85496 83648 86296 83768
rect 0 82968 800 83088
rect 85496 82288 86296 82408
rect 0 81608 800 81728
rect 85496 81608 86296 81728
rect 0 80248 800 80368
rect 85496 80248 86296 80368
rect 0 79568 800 79688
rect 85496 78888 86296 79008
rect 0 78208 800 78328
rect 85496 77528 86296 77648
rect 0 76848 800 76968
rect 85496 76168 86296 76288
rect 0 75488 800 75608
rect 85496 75488 86296 75608
rect 0 74128 800 74248
rect 85496 74128 86296 74248
rect 0 73448 800 73568
rect 85496 72768 86296 72888
rect 0 72088 800 72208
rect 85496 71408 86296 71528
rect 0 70728 800 70848
rect 85496 70048 86296 70168
rect 0 69368 800 69488
rect 85496 69368 86296 69488
rect 0 68008 800 68128
rect 85496 68008 86296 68128
rect 0 67328 800 67448
rect 85496 66648 86296 66768
rect 0 65968 800 66088
rect 85496 65288 86296 65408
rect 0 64608 800 64728
rect 85496 63928 86296 64048
rect 0 63248 800 63368
rect 85496 63248 86296 63368
rect 0 61888 800 62008
rect 85496 61888 86296 62008
rect 0 61208 800 61328
rect 85496 60528 86296 60648
rect 0 59848 800 59968
rect 85496 59168 86296 59288
rect 0 58488 800 58608
rect 85496 57808 86296 57928
rect 0 57128 800 57248
rect 85496 57128 86296 57248
rect 0 55768 800 55888
rect 85496 55768 86296 55888
rect 0 55088 800 55208
rect 85496 54408 86296 54528
rect 0 53728 800 53848
rect 85496 53048 86296 53168
rect 0 52368 800 52488
rect 85496 51688 86296 51808
rect 0 51008 800 51128
rect 85496 51008 86296 51128
rect 0 49648 800 49768
rect 85496 49648 86296 49768
rect 0 48968 800 49088
rect 85496 48288 86296 48408
rect 0 47608 800 47728
rect 85496 46928 86296 47048
rect 0 46248 800 46368
rect 85496 45568 86296 45688
rect 0 44888 800 45008
rect 85496 44888 86296 45008
rect 0 43528 800 43648
rect 85496 43528 86296 43648
rect 0 42848 800 42968
rect 85496 42168 86296 42288
rect 0 41488 800 41608
rect 85496 40808 86296 40928
rect 0 40128 800 40248
rect 85496 39448 86296 39568
rect 0 38768 800 38888
rect 85496 38768 86296 38888
rect 0 37408 800 37528
rect 85496 37408 86296 37528
rect 0 36728 800 36848
rect 85496 36048 86296 36168
rect 0 35368 800 35488
rect 85496 34688 86296 34808
rect 0 34008 800 34128
rect 85496 33328 86296 33448
rect 0 32648 800 32768
rect 85496 32648 86296 32768
rect 0 31288 800 31408
rect 85496 31288 86296 31408
rect 0 30608 800 30728
rect 85496 29928 86296 30048
rect 0 29248 800 29368
rect 85496 28568 86296 28688
rect 0 27888 800 28008
rect 85496 27208 86296 27328
rect 0 26528 800 26648
rect 85496 25848 86296 25968
rect 0 25168 800 25288
rect 85496 25168 86296 25288
rect 0 24488 800 24608
rect 85496 23808 86296 23928
rect 0 23128 800 23248
rect 85496 22448 86296 22568
rect 0 21768 800 21888
rect 85496 21088 86296 21208
rect 0 20408 800 20528
rect 85496 19728 86296 19848
rect 0 19048 800 19168
rect 85496 19048 86296 19168
rect 0 18368 800 18488
rect 85496 17688 86296 17808
rect 0 17008 800 17128
rect 85496 16328 86296 16448
rect 0 15648 800 15768
rect 85496 14968 86296 15088
rect 0 14288 800 14408
rect 85496 13608 86296 13728
rect 0 12928 800 13048
rect 85496 12928 86296 13048
rect 0 12248 800 12368
rect 85496 11568 86296 11688
rect 0 10888 800 11008
rect 85496 10208 86296 10328
rect 0 9528 800 9648
rect 85496 8848 86296 8968
rect 0 8168 800 8288
rect 85496 7488 86296 7608
rect 0 6808 800 6928
rect 85496 6808 86296 6928
rect 0 6128 800 6248
rect 85496 5448 86296 5568
rect 0 4768 800 4888
rect 85496 4088 86296 4208
rect 0 3408 800 3528
rect 85496 2728 86296 2848
rect 0 2048 800 2168
rect 85496 1368 86296 1488
rect 0 688 800 808
rect 85496 688 86296 808
<< obsm3 >>
rect 880 87648 85416 87821
rect 800 86568 85639 87648
rect 880 86288 85416 86568
rect 800 85888 85639 86288
rect 880 85608 85639 85888
rect 800 85208 85639 85608
rect 800 84928 85416 85208
rect 800 84528 85639 84928
rect 880 84248 85639 84528
rect 800 83848 85639 84248
rect 800 83568 85416 83848
rect 800 83168 85639 83568
rect 880 82888 85639 83168
rect 800 82488 85639 82888
rect 800 82208 85416 82488
rect 800 81808 85639 82208
rect 880 81528 85416 81808
rect 800 80448 85639 81528
rect 880 80168 85416 80448
rect 800 79768 85639 80168
rect 880 79488 85639 79768
rect 800 79088 85639 79488
rect 800 78808 85416 79088
rect 800 78408 85639 78808
rect 880 78128 85639 78408
rect 800 77728 85639 78128
rect 800 77448 85416 77728
rect 800 77048 85639 77448
rect 880 76768 85639 77048
rect 800 76368 85639 76768
rect 800 76088 85416 76368
rect 800 75688 85639 76088
rect 880 75408 85416 75688
rect 800 74328 85639 75408
rect 880 74048 85416 74328
rect 800 73648 85639 74048
rect 880 73368 85639 73648
rect 800 72968 85639 73368
rect 800 72688 85416 72968
rect 800 72288 85639 72688
rect 880 72008 85639 72288
rect 800 71608 85639 72008
rect 800 71328 85416 71608
rect 800 70928 85639 71328
rect 880 70648 85639 70928
rect 800 70248 85639 70648
rect 800 69968 85416 70248
rect 800 69568 85639 69968
rect 880 69288 85416 69568
rect 800 68208 85639 69288
rect 880 67928 85416 68208
rect 800 67528 85639 67928
rect 880 67248 85639 67528
rect 800 66848 85639 67248
rect 800 66568 85416 66848
rect 800 66168 85639 66568
rect 880 65888 85639 66168
rect 800 65488 85639 65888
rect 800 65208 85416 65488
rect 800 64808 85639 65208
rect 880 64528 85639 64808
rect 800 64128 85639 64528
rect 800 63848 85416 64128
rect 800 63448 85639 63848
rect 880 63168 85416 63448
rect 800 62088 85639 63168
rect 880 61808 85416 62088
rect 800 61408 85639 61808
rect 880 61128 85639 61408
rect 800 60728 85639 61128
rect 800 60448 85416 60728
rect 800 60048 85639 60448
rect 880 59768 85639 60048
rect 800 59368 85639 59768
rect 800 59088 85416 59368
rect 800 58688 85639 59088
rect 880 58408 85639 58688
rect 800 58008 85639 58408
rect 800 57728 85416 58008
rect 800 57328 85639 57728
rect 880 57048 85416 57328
rect 800 55968 85639 57048
rect 880 55688 85416 55968
rect 800 55288 85639 55688
rect 880 55008 85639 55288
rect 800 54608 85639 55008
rect 800 54328 85416 54608
rect 800 53928 85639 54328
rect 880 53648 85639 53928
rect 800 53248 85639 53648
rect 800 52968 85416 53248
rect 800 52568 85639 52968
rect 880 52288 85639 52568
rect 800 51888 85639 52288
rect 800 51608 85416 51888
rect 800 51208 85639 51608
rect 880 50928 85416 51208
rect 800 49848 85639 50928
rect 880 49568 85416 49848
rect 800 49168 85639 49568
rect 880 48888 85639 49168
rect 800 48488 85639 48888
rect 800 48208 85416 48488
rect 800 47808 85639 48208
rect 880 47528 85639 47808
rect 800 47128 85639 47528
rect 800 46848 85416 47128
rect 800 46448 85639 46848
rect 880 46168 85639 46448
rect 800 45768 85639 46168
rect 800 45488 85416 45768
rect 800 45088 85639 45488
rect 880 44808 85416 45088
rect 800 43728 85639 44808
rect 880 43448 85416 43728
rect 800 43048 85639 43448
rect 880 42768 85639 43048
rect 800 42368 85639 42768
rect 800 42088 85416 42368
rect 800 41688 85639 42088
rect 880 41408 85639 41688
rect 800 41008 85639 41408
rect 800 40728 85416 41008
rect 800 40328 85639 40728
rect 880 40048 85639 40328
rect 800 39648 85639 40048
rect 800 39368 85416 39648
rect 800 38968 85639 39368
rect 880 38688 85416 38968
rect 800 37608 85639 38688
rect 880 37328 85416 37608
rect 800 36928 85639 37328
rect 880 36648 85639 36928
rect 800 36248 85639 36648
rect 800 35968 85416 36248
rect 800 35568 85639 35968
rect 880 35288 85639 35568
rect 800 34888 85639 35288
rect 800 34608 85416 34888
rect 800 34208 85639 34608
rect 880 33928 85639 34208
rect 800 33528 85639 33928
rect 800 33248 85416 33528
rect 800 32848 85639 33248
rect 880 32568 85416 32848
rect 800 31488 85639 32568
rect 880 31208 85416 31488
rect 800 30808 85639 31208
rect 880 30528 85639 30808
rect 800 30128 85639 30528
rect 800 29848 85416 30128
rect 800 29448 85639 29848
rect 880 29168 85639 29448
rect 800 28768 85639 29168
rect 800 28488 85416 28768
rect 800 28088 85639 28488
rect 880 27808 85639 28088
rect 800 27408 85639 27808
rect 800 27128 85416 27408
rect 800 26728 85639 27128
rect 880 26448 85639 26728
rect 800 26048 85639 26448
rect 800 25768 85416 26048
rect 800 25368 85639 25768
rect 880 25088 85416 25368
rect 800 24688 85639 25088
rect 880 24408 85639 24688
rect 800 24008 85639 24408
rect 800 23728 85416 24008
rect 800 23328 85639 23728
rect 880 23048 85639 23328
rect 800 22648 85639 23048
rect 800 22368 85416 22648
rect 800 21968 85639 22368
rect 880 21688 85639 21968
rect 800 21288 85639 21688
rect 800 21008 85416 21288
rect 800 20608 85639 21008
rect 880 20328 85639 20608
rect 800 19928 85639 20328
rect 800 19648 85416 19928
rect 800 19248 85639 19648
rect 880 18968 85416 19248
rect 800 18568 85639 18968
rect 880 18288 85639 18568
rect 800 17888 85639 18288
rect 800 17608 85416 17888
rect 800 17208 85639 17608
rect 880 16928 85639 17208
rect 800 16528 85639 16928
rect 800 16248 85416 16528
rect 800 15848 85639 16248
rect 880 15568 85639 15848
rect 800 15168 85639 15568
rect 800 14888 85416 15168
rect 800 14488 85639 14888
rect 880 14208 85639 14488
rect 800 13808 85639 14208
rect 800 13528 85416 13808
rect 800 13128 85639 13528
rect 880 12848 85416 13128
rect 800 12448 85639 12848
rect 880 12168 85639 12448
rect 800 11768 85639 12168
rect 800 11488 85416 11768
rect 800 11088 85639 11488
rect 880 10808 85639 11088
rect 800 10408 85639 10808
rect 800 10128 85416 10408
rect 800 9728 85639 10128
rect 880 9448 85639 9728
rect 800 9048 85639 9448
rect 800 8768 85416 9048
rect 800 8368 85639 8768
rect 880 8088 85639 8368
rect 800 7688 85639 8088
rect 800 7408 85416 7688
rect 800 7008 85639 7408
rect 880 6728 85416 7008
rect 800 6328 85639 6728
rect 880 6048 85639 6328
rect 800 5648 85639 6048
rect 800 5368 85416 5648
rect 800 4968 85639 5368
rect 880 4688 85639 4968
rect 800 4288 85639 4688
rect 800 4008 85416 4288
rect 800 3608 85639 4008
rect 880 3328 85639 3608
rect 800 2928 85639 3328
rect 800 2648 85416 2928
rect 800 2248 85639 2648
rect 880 1968 85639 2248
rect 800 1568 85639 1968
rect 800 1288 85416 1568
rect 800 888 85639 1288
rect 880 715 85416 888
<< metal4 >>
rect 4208 2128 4528 86000
rect 4868 2128 5188 86000
rect 34928 2128 35248 86000
rect 35588 2128 35908 86000
rect 65648 2128 65968 86000
rect 66308 2128 66628 86000
<< obsm4 >>
rect 6683 86080 83845 86325
rect 6683 2048 34848 86080
rect 35328 2048 35508 86080
rect 35988 2048 65568 86080
rect 66048 2048 66228 86080
rect 66708 2048 83845 86080
rect 6683 1939 83845 2048
<< metal5 >>
rect 1056 67278 85240 67598
rect 1056 66618 85240 66938
rect 1056 36642 85240 36962
rect 1056 35982 85240 36302
rect 1056 6006 85240 6326
rect 1056 5346 85240 5666
<< obsm5 >>
rect 22748 23980 36316 24300
<< labels >>
rlabel metal4 s 4868 2128 5188 86000 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 86000 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 86000 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 85240 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 85240 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67278 85240 67598 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 86000 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 86000 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 86000 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 85240 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 85240 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 85240 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 30608 800 30728 6 clk
port 3 nsew signal input
rlabel metal3 s 85496 51008 86296 51128 6 cracked
port 4 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 done
port 5 nsew signal output
rlabel metal3 s 85496 60528 86296 60648 6 hash[0]
port 6 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 hash[100]
port 7 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 hash[101]
port 8 nsew signal input
rlabel metal2 s 23846 87640 23902 88440 6 hash[102]
port 9 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 hash[103]
port 10 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 hash[104]
port 11 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 hash[105]
port 12 nsew signal input
rlabel metal3 s 85496 49648 86296 49768 6 hash[106]
port 13 nsew signal input
rlabel metal2 s 16762 87640 16818 88440 6 hash[107]
port 14 nsew signal input
rlabel metal2 s 13542 87640 13598 88440 6 hash[108]
port 15 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 hash[109]
port 16 nsew signal input
rlabel metal2 s 43810 87640 43866 88440 6 hash[10]
port 17 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 hash[110]
port 18 nsew signal input
rlabel metal3 s 85496 37408 86296 37528 6 hash[111]
port 19 nsew signal input
rlabel metal2 s 64418 87640 64474 88440 6 hash[112]
port 20 nsew signal input
rlabel metal3 s 85496 51688 86296 51808 6 hash[113]
port 21 nsew signal input
rlabel metal2 s 20626 87640 20682 88440 6 hash[114]
port 22 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 hash[115]
port 23 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 hash[116]
port 24 nsew signal input
rlabel metal3 s 85496 55768 86296 55888 6 hash[117]
port 25 nsew signal input
rlabel metal3 s 85496 32648 86296 32768 6 hash[118]
port 26 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 hash[119]
port 27 nsew signal input
rlabel metal2 s 81806 87640 81862 88440 6 hash[11]
port 28 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 hash[120]
port 29 nsew signal input
rlabel metal2 s 14830 87640 14886 88440 6 hash[121]
port 30 nsew signal input
rlabel metal2 s 1950 87640 2006 88440 6 hash[122]
port 31 nsew signal input
rlabel metal2 s 52826 87640 52882 88440 6 hash[123]
port 32 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 hash[124]
port 33 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 hash[125]
port 34 nsew signal input
rlabel metal3 s 85496 4088 86296 4208 6 hash[126]
port 35 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 hash[127]
port 36 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 hash[128]
port 37 nsew signal input
rlabel metal3 s 85496 61888 86296 62008 6 hash[129]
port 38 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 hash[12]
port 39 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 hash[130]
port 40 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 hash[131]
port 41 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 hash[132]
port 42 nsew signal input
rlabel metal3 s 85496 82288 86296 82408 6 hash[133]
port 43 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 hash[134]
port 44 nsew signal input
rlabel metal3 s 0 688 800 808 6 hash[135]
port 45 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 hash[136]
port 46 nsew signal input
rlabel metal2 s 7746 87640 7802 88440 6 hash[137]
port 47 nsew signal input
rlabel metal3 s 85496 76168 86296 76288 6 hash[138]
port 48 nsew signal input
rlabel metal2 s 33506 87640 33562 88440 6 hash[139]
port 49 nsew signal input
rlabel metal2 s 42522 87640 42578 88440 6 hash[13]
port 50 nsew signal input
rlabel metal3 s 85496 78888 86296 79008 6 hash[140]
port 51 nsew signal input
rlabel metal2 s 19338 87640 19394 88440 6 hash[141]
port 52 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 hash[142]
port 53 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 hash[143]
port 54 nsew signal input
rlabel metal2 s 41234 87640 41290 88440 6 hash[144]
port 55 nsew signal input
rlabel metal3 s 85496 1368 86296 1488 6 hash[145]
port 56 nsew signal input
rlabel metal3 s 85496 86368 86296 86488 6 hash[146]
port 57 nsew signal input
rlabel metal3 s 85496 38768 86296 38888 6 hash[147]
port 58 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 hash[148]
port 59 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 hash[149]
port 60 nsew signal input
rlabel metal2 s 55402 87640 55458 88440 6 hash[14]
port 61 nsew signal input
rlabel metal3 s 85496 69368 86296 69488 6 hash[150]
port 62 nsew signal input
rlabel metal3 s 85496 57128 86296 57248 6 hash[151]
port 63 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 hash[152]
port 64 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 hash[153]
port 65 nsew signal input
rlabel metal2 s 32218 87640 32274 88440 6 hash[154]
port 66 nsew signal input
rlabel metal2 s 27066 87640 27122 88440 6 hash[155]
port 67 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 hash[156]
port 68 nsew signal input
rlabel metal3 s 85496 70048 86296 70168 6 hash[157]
port 69 nsew signal input
rlabel metal3 s 85496 17688 86296 17808 6 hash[158]
port 70 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 hash[159]
port 71 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 hash[15]
port 72 nsew signal input
rlabel metal3 s 85496 10208 86296 10328 6 hash[160]
port 73 nsew signal input
rlabel metal3 s 85496 83648 86296 83768 6 hash[161]
port 74 nsew signal input
rlabel metal2 s 3238 87640 3294 88440 6 hash[162]
port 75 nsew signal input
rlabel metal3 s 85496 13608 86296 13728 6 hash[163]
port 76 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 hash[164]
port 77 nsew signal input
rlabel metal2 s 66994 87640 67050 88440 6 hash[165]
port 78 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 hash[166]
port 79 nsew signal input
rlabel metal2 s 21270 87640 21326 88440 6 hash[167]
port 80 nsew signal input
rlabel metal2 s 36726 87640 36782 88440 6 hash[168]
port 81 nsew signal input
rlabel metal3 s 85496 46928 86296 47048 6 hash[169]
port 82 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 hash[16]
port 83 nsew signal input
rlabel metal3 s 85496 14968 86296 15088 6 hash[170]
port 84 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 hash[171]
port 85 nsew signal input
rlabel metal2 s 74722 87640 74778 88440 6 hash[172]
port 86 nsew signal input
rlabel metal2 s 28354 87640 28410 88440 6 hash[173]
port 87 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 hash[174]
port 88 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 hash[175]
port 89 nsew signal input
rlabel metal3 s 85496 75488 86296 75608 6 hash[176]
port 90 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 hash[177]
port 91 nsew signal input
rlabel metal3 s 85496 25168 86296 25288 6 hash[178]
port 92 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 hash[179]
port 93 nsew signal input
rlabel metal2 s 29642 87640 29698 88440 6 hash[17]
port 94 nsew signal input
rlabel metal3 s 85496 25848 86296 25968 6 hash[180]
port 95 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 hash[181]
port 96 nsew signal input
rlabel metal3 s 85496 27208 86296 27328 6 hash[182]
port 97 nsew signal input
rlabel metal2 s 39946 87640 40002 88440 6 hash[183]
port 98 nsew signal input
rlabel metal2 s 85670 87640 85726 88440 6 hash[184]
port 99 nsew signal input
rlabel metal3 s 85496 77528 86296 77648 6 hash[185]
port 100 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 hash[186]
port 101 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 hash[187]
port 102 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 hash[188]
port 103 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 hash[189]
port 104 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 hash[18]
port 105 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 hash[190]
port 106 nsew signal input
rlabel metal2 s 18050 87640 18106 88440 6 hash[191]
port 107 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 hash[192]
port 108 nsew signal input
rlabel metal2 s 80518 87640 80574 88440 6 hash[193]
port 109 nsew signal input
rlabel metal3 s 85496 2728 86296 2848 6 hash[194]
port 110 nsew signal input
rlabel metal3 s 85496 59168 86296 59288 6 hash[195]
port 111 nsew signal input
rlabel metal3 s 85496 22448 86296 22568 6 hash[196]
port 112 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 hash[197]
port 113 nsew signal input
rlabel metal2 s 45098 87640 45154 88440 6 hash[198]
port 114 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 hash[199]
port 115 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 hash[19]
port 116 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 hash[1]
port 117 nsew signal input
rlabel metal2 s 78586 87640 78642 88440 6 hash[200]
port 118 nsew signal input
rlabel metal2 s 26422 87640 26478 88440 6 hash[201]
port 119 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 hash[202]
port 120 nsew signal input
rlabel metal3 s 85496 688 86296 808 6 hash[203]
port 121 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 hash[204]
port 122 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 hash[205]
port 123 nsew signal input
rlabel metal3 s 85496 68008 86296 68128 6 hash[206]
port 124 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 hash[207]
port 125 nsew signal input
rlabel metal3 s 85496 8848 86296 8968 6 hash[208]
port 126 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 hash[209]
port 127 nsew signal input
rlabel metal2 s 65706 87640 65762 88440 6 hash[20]
port 128 nsew signal input
rlabel metal2 s 51538 87640 51594 88440 6 hash[210]
port 129 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 hash[211]
port 130 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 hash[212]
port 131 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 hash[213]
port 132 nsew signal input
rlabel metal3 s 85496 7488 86296 7608 6 hash[214]
port 133 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 hash[215]
port 134 nsew signal input
rlabel metal3 s 85496 48288 86296 48408 6 hash[216]
port 135 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 hash[217]
port 136 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 hash[218]
port 137 nsew signal input
rlabel metal2 s 68282 87640 68338 88440 6 hash[219]
port 138 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 hash[21]
port 139 nsew signal input
rlabel metal2 s 72790 87640 72846 88440 6 hash[220]
port 140 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 hash[221]
port 141 nsew signal input
rlabel metal3 s 85496 11568 86296 11688 6 hash[222]
port 142 nsew signal input
rlabel metal3 s 85496 40808 86296 40928 6 hash[223]
port 143 nsew signal input
rlabel metal3 s 85496 45568 86296 45688 6 hash[224]
port 144 nsew signal input
rlabel metal2 s 12254 87640 12310 88440 6 hash[225]
port 145 nsew signal input
rlabel metal3 s 85496 85008 86296 85128 6 hash[226]
port 146 nsew signal input
rlabel metal2 s 48318 87640 48374 88440 6 hash[227]
port 147 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 hash[228]
port 148 nsew signal input
rlabel metal3 s 85496 54408 86296 54528 6 hash[229]
port 149 nsew signal input
rlabel metal2 s 76010 87640 76066 88440 6 hash[22]
port 150 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 hash[230]
port 151 nsew signal input
rlabel metal2 s 34150 87640 34206 88440 6 hash[231]
port 152 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 hash[232]
port 153 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 hash[233]
port 154 nsew signal input
rlabel metal3 s 85496 53048 86296 53168 6 hash[234]
port 155 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 hash[235]
port 156 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 hash[236]
port 157 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 hash[237]
port 158 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 hash[238]
port 159 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 hash[239]
port 160 nsew signal input
rlabel metal3 s 85496 63928 86296 64048 6 hash[23]
port 161 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 hash[240]
port 162 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 hash[241]
port 163 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 hash[242]
port 164 nsew signal input
rlabel metal3 s 85496 16328 86296 16448 6 hash[243]
port 165 nsew signal input
rlabel metal3 s 85496 29928 86296 30048 6 hash[244]
port 166 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 hash[245]
port 167 nsew signal input
rlabel metal2 s 70214 87640 70270 88440 6 hash[246]
port 168 nsew signal input
rlabel metal2 s 45742 87640 45798 88440 6 hash[247]
port 169 nsew signal input
rlabel metal3 s 85496 28568 86296 28688 6 hash[248]
port 170 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 hash[249]
port 171 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 hash[24]
port 172 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 hash[250]
port 173 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 hash[251]
port 174 nsew signal input
rlabel metal2 s 662 87640 718 88440 6 hash[252]
port 175 nsew signal input
rlabel metal2 s 9034 87640 9090 88440 6 hash[253]
port 176 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 hash[254]
port 177 nsew signal input
rlabel metal2 s 59910 87640 59966 88440 6 hash[255]
port 178 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 hash[25]
port 179 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 hash[26]
port 180 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 hash[27]
port 181 nsew signal input
rlabel metal3 s 85496 33328 86296 33448 6 hash[28]
port 182 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 hash[29]
port 183 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 hash[2]
port 184 nsew signal input
rlabel metal2 s 61198 87640 61254 88440 6 hash[30]
port 185 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 hash[31]
port 186 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 hash[32]
port 187 nsew signal input
rlabel metal2 s 56690 87640 56746 88440 6 hash[33]
port 188 nsew signal input
rlabel metal2 s 62486 87640 62542 88440 6 hash[34]
port 189 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 hash[35]
port 190 nsew signal input
rlabel metal2 s 50894 87640 50950 88440 6 hash[36]
port 191 nsew signal input
rlabel metal2 s 25134 87640 25190 88440 6 hash[37]
port 192 nsew signal input
rlabel metal2 s 5170 87640 5226 88440 6 hash[38]
port 193 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 hash[39]
port 194 nsew signal input
rlabel metal2 s 39302 87640 39358 88440 6 hash[3]
port 195 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 hash[40]
port 196 nsew signal input
rlabel metal2 s 15474 87640 15530 88440 6 hash[41]
port 197 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 hash[42]
port 198 nsew signal input
rlabel metal3 s 85496 39448 86296 39568 6 hash[43]
port 199 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 hash[44]
port 200 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 hash[45]
port 201 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 hash[46]
port 202 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 hash[47]
port 203 nsew signal input
rlabel metal2 s 79874 87640 79930 88440 6 hash[48]
port 204 nsew signal input
rlabel metal3 s 85496 72768 86296 72888 6 hash[49]
port 205 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 hash[4]
port 206 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 hash[50]
port 207 nsew signal input
rlabel metal3 s 85496 6808 86296 6928 6 hash[51]
port 208 nsew signal input
rlabel metal2 s 38014 87640 38070 88440 6 hash[52]
port 209 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 hash[53]
port 210 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 hash[54]
port 211 nsew signal input
rlabel metal2 s 54114 87640 54170 88440 6 hash[55]
port 212 nsew signal input
rlabel metal3 s 85496 36048 86296 36168 6 hash[56]
port 213 nsew signal input
rlabel metal3 s 85496 66648 86296 66768 6 hash[57]
port 214 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 hash[58]
port 215 nsew signal input
rlabel metal3 s 85496 87728 86296 87848 6 hash[59]
port 216 nsew signal input
rlabel metal3 s 85496 23808 86296 23928 6 hash[5]
port 217 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 hash[60]
port 218 nsew signal input
rlabel metal2 s 84382 87640 84438 88440 6 hash[61]
port 219 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 hash[62]
port 220 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 hash[63]
port 221 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 hash[64]
port 222 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 hash[65]
port 223 nsew signal input
rlabel metal3 s 85496 12928 86296 13048 6 hash[66]
port 224 nsew signal input
rlabel metal2 s 47030 87640 47086 88440 6 hash[67]
port 225 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 hash[68]
port 226 nsew signal input
rlabel metal2 s 3882 87640 3938 88440 6 hash[69]
port 227 nsew signal input
rlabel metal2 s 9678 87640 9734 88440 6 hash[6]
port 228 nsew signal input
rlabel metal2 s 6458 87640 6514 88440 6 hash[70]
port 229 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 hash[71]
port 230 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 hash[72]
port 231 nsew signal input
rlabel metal3 s 85496 34688 86296 34808 6 hash[73]
port 232 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 hash[74]
port 233 nsew signal input
rlabel metal2 s 74078 87640 74134 88440 6 hash[75]
port 234 nsew signal input
rlabel metal3 s 85496 81608 86296 81728 6 hash[76]
port 235 nsew signal input
rlabel metal2 s 22558 87640 22614 88440 6 hash[77]
port 236 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 hash[78]
port 237 nsew signal input
rlabel metal3 s 85496 43528 86296 43648 6 hash[79]
port 238 nsew signal input
rlabel metal3 s 85496 80248 86296 80368 6 hash[7]
port 239 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 hash[80]
port 240 nsew signal input
rlabel metal3 s 85496 57808 86296 57928 6 hash[81]
port 241 nsew signal input
rlabel metal3 s 85496 19728 86296 19848 6 hash[82]
port 242 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 hash[83]
port 243 nsew signal input
rlabel metal2 s 83094 87640 83150 88440 6 hash[84]
port 244 nsew signal input
rlabel metal2 s 35438 87640 35494 88440 6 hash[85]
port 245 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 hash[86]
port 246 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 hash[87]
port 247 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 hash[88]
port 248 nsew signal input
rlabel metal3 s 85496 19048 86296 19168 6 hash[89]
port 249 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 hash[8]
port 250 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 hash[90]
port 251 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 hash[91]
port 252 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 hash[92]
port 253 nsew signal input
rlabel metal3 s 85496 31288 86296 31408 6 hash[93]
port 254 nsew signal input
rlabel metal2 s 77298 87640 77354 88440 6 hash[94]
port 255 nsew signal input
rlabel metal3 s 85496 71408 86296 71528 6 hash[95]
port 256 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 hash[96]
port 257 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 hash[97]
port 258 nsew signal input
rlabel metal3 s 85496 44888 86296 45008 6 hash[98]
port 259 nsew signal input
rlabel metal2 s 662 0 718 800 6 hash[99]
port 260 nsew signal input
rlabel metal3 s 85496 74128 86296 74248 6 hash[9]
port 261 nsew signal input
rlabel metal2 s 71502 87640 71558 88440 6 init
port 262 nsew signal input
rlabel metal3 s 85496 5448 86296 5568 6 password_count[0]
port 263 nsew signal output
rlabel metal2 s 68926 87640 68982 88440 6 password_count[10]
port 264 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 password_count[11]
port 265 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 password_count[12]
port 266 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 password_count[13]
port 267 nsew signal output
rlabel metal2 s 18 0 74 800 6 password_count[14]
port 268 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 password_count[15]
port 269 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 password_count[16]
port 270 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 password_count[17]
port 271 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 password_count[18]
port 272 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 password_count[19]
port 273 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 password_count[1]
port 274 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 password_count[20]
port 275 nsew signal output
rlabel metal2 s 49606 87640 49662 88440 6 password_count[21]
port 276 nsew signal output
rlabel metal2 s 30930 87640 30986 88440 6 password_count[22]
port 277 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 password_count[23]
port 278 nsew signal output
rlabel metal2 s 63130 87640 63186 88440 6 password_count[24]
port 279 nsew signal output
rlabel metal3 s 85496 21088 86296 21208 6 password_count[25]
port 280 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 password_count[26]
port 281 nsew signal output
rlabel metal3 s 85496 65288 86296 65408 6 password_count[27]
port 282 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 password_count[28]
port 283 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 password_count[29]
port 284 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 password_count[2]
port 285 nsew signal output
rlabel metal3 s 85496 63248 86296 63368 6 password_count[30]
port 286 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 password_count[31]
port 287 nsew signal output
rlabel metal2 s 58622 87640 58678 88440 6 password_count[3]
port 288 nsew signal output
rlabel metal2 s 57334 87640 57390 88440 6 password_count[4]
port 289 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 password_count[5]
port 290 nsew signal output
rlabel metal2 s 10966 87640 11022 88440 6 password_count[6]
port 291 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 password_count[7]
port 292 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 password_count[8]
port 293 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 password_count[9]
port 294 nsew signal output
rlabel metal3 s 85496 42168 86296 42288 6 reset
port 295 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 86296 88440
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 21864868
string GDS_FILE /openlane/designs/password_cracker/runs/RUN_2023.03.23_09.07.37/results/signoff/password_cracker.magic.gds
string GDS_START 944678
<< end >>

