VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO password_cracker
  CLASS BLOCK ;
  FOREIGN password_cracker ;
  ORIGIN 0.000 0.000 ;
  SIZE 431.480 BY 442.200 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 430.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 430.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 430.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 426.200 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 426.200 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 426.200 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 430.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 430.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 430.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 426.200 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 426.200 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 426.200 334.690 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END clk
  PIN cracked
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 255.040 431.480 255.640 ;
    END
  END cracked
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END done
  PIN hash[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 302.640 431.480 303.240 ;
    END
  END hash[0]
  PIN hash[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END hash[100]
  PIN hash[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END hash[101]
  PIN hash[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 438.200 119.510 442.200 ;
    END
  END hash[102]
  PIN hash[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END hash[103]
  PIN hash[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END hash[104]
  PIN hash[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END hash[105]
  PIN hash[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 248.240 431.480 248.840 ;
    END
  END hash[106]
  PIN hash[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 438.200 84.090 442.200 ;
    END
  END hash[107]
  PIN hash[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 438.200 67.990 442.200 ;
    END
  END hash[108]
  PIN hash[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END hash[109]
  PIN hash[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 438.200 219.330 442.200 ;
    END
  END hash[10]
  PIN hash[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END hash[110]
  PIN hash[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 187.040 431.480 187.640 ;
    END
  END hash[111]
  PIN hash[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 438.200 322.370 442.200 ;
    END
  END hash[112]
  PIN hash[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 258.440 431.480 259.040 ;
    END
  END hash[113]
  PIN hash[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 438.200 103.410 442.200 ;
    END
  END hash[114]
  PIN hash[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END hash[115]
  PIN hash[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END hash[116]
  PIN hash[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 278.840 431.480 279.440 ;
    END
  END hash[117]
  PIN hash[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 163.240 431.480 163.840 ;
    END
  END hash[118]
  PIN hash[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END hash[119]
  PIN hash[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 438.200 409.310 442.200 ;
    END
  END hash[11]
  PIN hash[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END hash[120]
  PIN hash[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 438.200 74.430 442.200 ;
    END
  END hash[121]
  PIN hash[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 438.200 10.030 442.200 ;
    END
  END hash[122]
  PIN hash[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 438.200 264.410 442.200 ;
    END
  END hash[123]
  PIN hash[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END hash[124]
  PIN hash[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END hash[125]
  PIN hash[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 20.440 431.480 21.040 ;
    END
  END hash[126]
  PIN hash[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END hash[127]
  PIN hash[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END hash[128]
  PIN hash[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 309.440 431.480 310.040 ;
    END
  END hash[129]
  PIN hash[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END hash[12]
  PIN hash[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END hash[130]
  PIN hash[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END hash[131]
  PIN hash[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END hash[132]
  PIN hash[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 411.440 431.480 412.040 ;
    END
  END hash[133]
  PIN hash[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END hash[134]
  PIN hash[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END hash[135]
  PIN hash[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END hash[136]
  PIN hash[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 438.200 39.010 442.200 ;
    END
  END hash[137]
  PIN hash[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 380.840 431.480 381.440 ;
    END
  END hash[138]
  PIN hash[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 438.200 167.810 442.200 ;
    END
  END hash[139]
  PIN hash[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 438.200 212.890 442.200 ;
    END
  END hash[13]
  PIN hash[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 394.440 431.480 395.040 ;
    END
  END hash[140]
  PIN hash[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 438.200 96.970 442.200 ;
    END
  END hash[141]
  PIN hash[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END hash[142]
  PIN hash[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END hash[143]
  PIN hash[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 438.200 206.450 442.200 ;
    END
  END hash[144]
  PIN hash[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 6.840 431.480 7.440 ;
    END
  END hash[145]
  PIN hash[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 431.840 431.480 432.440 ;
    END
  END hash[146]
  PIN hash[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 193.840 431.480 194.440 ;
    END
  END hash[147]
  PIN hash[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END hash[148]
  PIN hash[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END hash[149]
  PIN hash[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 438.200 277.290 442.200 ;
    END
  END hash[14]
  PIN hash[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 346.840 431.480 347.440 ;
    END
  END hash[150]
  PIN hash[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 285.640 431.480 286.240 ;
    END
  END hash[151]
  PIN hash[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END hash[152]
  PIN hash[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END hash[153]
  PIN hash[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 438.200 161.370 442.200 ;
    END
  END hash[154]
  PIN hash[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 438.200 135.610 442.200 ;
    END
  END hash[155]
  PIN hash[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END hash[156]
  PIN hash[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 350.240 431.480 350.840 ;
    END
  END hash[157]
  PIN hash[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 88.440 431.480 89.040 ;
    END
  END hash[158]
  PIN hash[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END hash[159]
  PIN hash[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END hash[15]
  PIN hash[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 51.040 431.480 51.640 ;
    END
  END hash[160]
  PIN hash[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 418.240 431.480 418.840 ;
    END
  END hash[161]
  PIN hash[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 438.200 16.470 442.200 ;
    END
  END hash[162]
  PIN hash[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 68.040 431.480 68.640 ;
    END
  END hash[163]
  PIN hash[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END hash[164]
  PIN hash[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 438.200 335.250 442.200 ;
    END
  END hash[165]
  PIN hash[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END hash[166]
  PIN hash[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 438.200 106.630 442.200 ;
    END
  END hash[167]
  PIN hash[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 438.200 183.910 442.200 ;
    END
  END hash[168]
  PIN hash[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 234.640 431.480 235.240 ;
    END
  END hash[169]
  PIN hash[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END hash[16]
  PIN hash[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 74.840 431.480 75.440 ;
    END
  END hash[170]
  PIN hash[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END hash[171]
  PIN hash[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 438.200 373.890 442.200 ;
    END
  END hash[172]
  PIN hash[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 438.200 142.050 442.200 ;
    END
  END hash[173]
  PIN hash[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END hash[174]
  PIN hash[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END hash[175]
  PIN hash[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 377.440 431.480 378.040 ;
    END
  END hash[176]
  PIN hash[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END hash[177]
  PIN hash[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 125.840 431.480 126.440 ;
    END
  END hash[178]
  PIN hash[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END hash[179]
  PIN hash[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 438.200 148.490 442.200 ;
    END
  END hash[17]
  PIN hash[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 129.240 431.480 129.840 ;
    END
  END hash[180]
  PIN hash[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END hash[181]
  PIN hash[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 136.040 431.480 136.640 ;
    END
  END hash[182]
  PIN hash[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 438.200 200.010 442.200 ;
    END
  END hash[183]
  PIN hash[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 438.200 428.630 442.200 ;
    END
  END hash[184]
  PIN hash[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 387.640 431.480 388.240 ;
    END
  END hash[185]
  PIN hash[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END hash[186]
  PIN hash[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END hash[187]
  PIN hash[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END hash[188]
  PIN hash[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END hash[189]
  PIN hash[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END hash[18]
  PIN hash[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END hash[190]
  PIN hash[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 438.200 90.530 442.200 ;
    END
  END hash[191]
  PIN hash[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END hash[192]
  PIN hash[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 438.200 402.870 442.200 ;
    END
  END hash[193]
  PIN hash[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 13.640 431.480 14.240 ;
    END
  END hash[194]
  PIN hash[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 295.840 431.480 296.440 ;
    END
  END hash[195]
  PIN hash[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 112.240 431.480 112.840 ;
    END
  END hash[196]
  PIN hash[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END hash[197]
  PIN hash[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 438.200 225.770 442.200 ;
    END
  END hash[198]
  PIN hash[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END hash[199]
  PIN hash[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END hash[19]
  PIN hash[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END hash[1]
  PIN hash[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 438.200 393.210 442.200 ;
    END
  END hash[200]
  PIN hash[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 438.200 132.390 442.200 ;
    END
  END hash[201]
  PIN hash[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END hash[202]
  PIN hash[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 3.440 431.480 4.040 ;
    END
  END hash[203]
  PIN hash[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END hash[204]
  PIN hash[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END hash[205]
  PIN hash[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 340.040 431.480 340.640 ;
    END
  END hash[206]
  PIN hash[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END hash[207]
  PIN hash[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 44.240 431.480 44.840 ;
    END
  END hash[208]
  PIN hash[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END hash[209]
  PIN hash[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 438.200 328.810 442.200 ;
    END
  END hash[20]
  PIN hash[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 438.200 257.970 442.200 ;
    END
  END hash[210]
  PIN hash[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END hash[211]
  PIN hash[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END hash[212]
  PIN hash[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END hash[213]
  PIN hash[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 37.440 431.480 38.040 ;
    END
  END hash[214]
  PIN hash[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END hash[215]
  PIN hash[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 241.440 431.480 242.040 ;
    END
  END hash[216]
  PIN hash[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END hash[217]
  PIN hash[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END hash[218]
  PIN hash[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 438.200 341.690 442.200 ;
    END
  END hash[219]
  PIN hash[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END hash[21]
  PIN hash[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 438.200 364.230 442.200 ;
    END
  END hash[220]
  PIN hash[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END hash[221]
  PIN hash[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 57.840 431.480 58.440 ;
    END
  END hash[222]
  PIN hash[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 204.040 431.480 204.640 ;
    END
  END hash[223]
  PIN hash[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 227.840 431.480 228.440 ;
    END
  END hash[224]
  PIN hash[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 438.200 61.550 442.200 ;
    END
  END hash[225]
  PIN hash[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 425.040 431.480 425.640 ;
    END
  END hash[226]
  PIN hash[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 438.200 241.870 442.200 ;
    END
  END hash[227]
  PIN hash[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END hash[228]
  PIN hash[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 272.040 431.480 272.640 ;
    END
  END hash[229]
  PIN hash[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 438.200 380.330 442.200 ;
    END
  END hash[22]
  PIN hash[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END hash[230]
  PIN hash[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 438.200 171.030 442.200 ;
    END
  END hash[231]
  PIN hash[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END hash[232]
  PIN hash[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END hash[233]
  PIN hash[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 265.240 431.480 265.840 ;
    END
  END hash[234]
  PIN hash[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END hash[235]
  PIN hash[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END hash[236]
  PIN hash[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END hash[237]
  PIN hash[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END hash[238]
  PIN hash[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END hash[239]
  PIN hash[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 319.640 431.480 320.240 ;
    END
  END hash[23]
  PIN hash[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END hash[240]
  PIN hash[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END hash[241]
  PIN hash[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END hash[242]
  PIN hash[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 81.640 431.480 82.240 ;
    END
  END hash[243]
  PIN hash[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 149.640 431.480 150.240 ;
    END
  END hash[244]
  PIN hash[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END hash[245]
  PIN hash[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 438.200 351.350 442.200 ;
    END
  END hash[246]
  PIN hash[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 438.200 228.990 442.200 ;
    END
  END hash[247]
  PIN hash[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 142.840 431.480 143.440 ;
    END
  END hash[248]
  PIN hash[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END hash[249]
  PIN hash[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END hash[24]
  PIN hash[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END hash[250]
  PIN hash[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END hash[251]
  PIN hash[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 438.200 3.590 442.200 ;
    END
  END hash[252]
  PIN hash[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 438.200 45.450 442.200 ;
    END
  END hash[253]
  PIN hash[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END hash[254]
  PIN hash[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 438.200 299.830 442.200 ;
    END
  END hash[255]
  PIN hash[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END hash[25]
  PIN hash[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END hash[26]
  PIN hash[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END hash[27]
  PIN hash[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 166.640 431.480 167.240 ;
    END
  END hash[28]
  PIN hash[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END hash[29]
  PIN hash[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END hash[2]
  PIN hash[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 438.200 306.270 442.200 ;
    END
  END hash[30]
  PIN hash[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END hash[31]
  PIN hash[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END hash[32]
  PIN hash[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 438.200 283.730 442.200 ;
    END
  END hash[33]
  PIN hash[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 438.200 312.710 442.200 ;
    END
  END hash[34]
  PIN hash[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END hash[35]
  PIN hash[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 438.200 254.750 442.200 ;
    END
  END hash[36]
  PIN hash[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 438.200 125.950 442.200 ;
    END
  END hash[37]
  PIN hash[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 438.200 26.130 442.200 ;
    END
  END hash[38]
  PIN hash[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END hash[39]
  PIN hash[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 438.200 196.790 442.200 ;
    END
  END hash[3]
  PIN hash[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END hash[40]
  PIN hash[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 438.200 77.650 442.200 ;
    END
  END hash[41]
  PIN hash[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END hash[42]
  PIN hash[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 197.240 431.480 197.840 ;
    END
  END hash[43]
  PIN hash[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END hash[44]
  PIN hash[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END hash[45]
  PIN hash[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END hash[46]
  PIN hash[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END hash[47]
  PIN hash[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 438.200 399.650 442.200 ;
    END
  END hash[48]
  PIN hash[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 363.840 431.480 364.440 ;
    END
  END hash[49]
  PIN hash[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END hash[4]
  PIN hash[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END hash[50]
  PIN hash[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 34.040 431.480 34.640 ;
    END
  END hash[51]
  PIN hash[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 438.200 190.350 442.200 ;
    END
  END hash[52]
  PIN hash[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END hash[53]
  PIN hash[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END hash[54]
  PIN hash[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 438.200 270.850 442.200 ;
    END
  END hash[55]
  PIN hash[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 180.240 431.480 180.840 ;
    END
  END hash[56]
  PIN hash[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 333.240 431.480 333.840 ;
    END
  END hash[57]
  PIN hash[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END hash[58]
  PIN hash[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 438.640 431.480 439.240 ;
    END
  END hash[59]
  PIN hash[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 119.040 431.480 119.640 ;
    END
  END hash[5]
  PIN hash[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END hash[60]
  PIN hash[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 438.200 422.190 442.200 ;
    END
  END hash[61]
  PIN hash[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END hash[62]
  PIN hash[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END hash[63]
  PIN hash[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END hash[64]
  PIN hash[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END hash[65]
  PIN hash[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 64.640 431.480 65.240 ;
    END
  END hash[66]
  PIN hash[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 438.200 235.430 442.200 ;
    END
  END hash[67]
  PIN hash[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END hash[68]
  PIN hash[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 438.200 19.690 442.200 ;
    END
  END hash[69]
  PIN hash[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 438.200 48.670 442.200 ;
    END
  END hash[6]
  PIN hash[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 438.200 32.570 442.200 ;
    END
  END hash[70]
  PIN hash[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END hash[71]
  PIN hash[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END hash[72]
  PIN hash[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 173.440 431.480 174.040 ;
    END
  END hash[73]
  PIN hash[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END hash[74]
  PIN hash[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 438.200 370.670 442.200 ;
    END
  END hash[75]
  PIN hash[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 408.040 431.480 408.640 ;
    END
  END hash[76]
  PIN hash[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 438.200 113.070 442.200 ;
    END
  END hash[77]
  PIN hash[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END hash[78]
  PIN hash[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 217.640 431.480 218.240 ;
    END
  END hash[79]
  PIN hash[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 401.240 431.480 401.840 ;
    END
  END hash[7]
  PIN hash[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END hash[80]
  PIN hash[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 289.040 431.480 289.640 ;
    END
  END hash[81]
  PIN hash[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 98.640 431.480 99.240 ;
    END
  END hash[82]
  PIN hash[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END hash[83]
  PIN hash[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 438.200 415.750 442.200 ;
    END
  END hash[84]
  PIN hash[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 438.200 177.470 442.200 ;
    END
  END hash[85]
  PIN hash[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END hash[86]
  PIN hash[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END hash[87]
  PIN hash[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END hash[88]
  PIN hash[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 95.240 431.480 95.840 ;
    END
  END hash[89]
  PIN hash[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END hash[8]
  PIN hash[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END hash[90]
  PIN hash[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END hash[91]
  PIN hash[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END hash[92]
  PIN hash[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 156.440 431.480 157.040 ;
    END
  END hash[93]
  PIN hash[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 438.200 386.770 442.200 ;
    END
  END hash[94]
  PIN hash[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 357.040 431.480 357.640 ;
    END
  END hash[95]
  PIN hash[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END hash[96]
  PIN hash[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END hash[97]
  PIN hash[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 224.440 431.480 225.040 ;
    END
  END hash[98]
  PIN hash[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END hash[99]
  PIN hash[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 370.640 431.480 371.240 ;
    END
  END hash[9]
  PIN init
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 438.200 357.790 442.200 ;
    END
  END init
  PIN password_count[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 27.240 431.480 27.840 ;
    END
  END password_count[0]
  PIN password_count[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 438.200 344.910 442.200 ;
    END
  END password_count[10]
  PIN password_count[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END password_count[11]
  PIN password_count[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END password_count[12]
  PIN password_count[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END password_count[13]
  PIN password_count[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END password_count[14]
  PIN password_count[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END password_count[15]
  PIN password_count[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END password_count[16]
  PIN password_count[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END password_count[17]
  PIN password_count[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END password_count[18]
  PIN password_count[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END password_count[19]
  PIN password_count[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END password_count[1]
  PIN password_count[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END password_count[20]
  PIN password_count[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 438.200 248.310 442.200 ;
    END
  END password_count[21]
  PIN password_count[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 438.200 154.930 442.200 ;
    END
  END password_count[22]
  PIN password_count[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END password_count[23]
  PIN password_count[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 438.200 315.930 442.200 ;
    END
  END password_count[24]
  PIN password_count[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 105.440 431.480 106.040 ;
    END
  END password_count[25]
  PIN password_count[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END password_count[26]
  PIN password_count[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 326.440 431.480 327.040 ;
    END
  END password_count[27]
  PIN password_count[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END password_count[28]
  PIN password_count[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END password_count[29]
  PIN password_count[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END password_count[2]
  PIN password_count[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 316.240 431.480 316.840 ;
    END
  END password_count[30]
  PIN password_count[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END password_count[31]
  PIN password_count[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 438.200 293.390 442.200 ;
    END
  END password_count[3]
  PIN password_count[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 438.200 286.950 442.200 ;
    END
  END password_count[4]
  PIN password_count[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END password_count[5]
  PIN password_count[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 438.200 55.110 442.200 ;
    END
  END password_count[6]
  PIN password_count[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END password_count[7]
  PIN password_count[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END password_count[8]
  PIN password_count[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END password_count[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.480 210.840 431.480 211.440 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 425.960 429.845 ;
      LAYER met1 ;
        RECT 0.070 7.860 430.490 437.200 ;
      LAYER met2 ;
        RECT 0.100 437.920 3.030 439.125 ;
        RECT 3.870 437.920 9.470 439.125 ;
        RECT 10.310 437.920 15.910 439.125 ;
        RECT 16.750 437.920 19.130 439.125 ;
        RECT 19.970 437.920 25.570 439.125 ;
        RECT 26.410 437.920 32.010 439.125 ;
        RECT 32.850 437.920 38.450 439.125 ;
        RECT 39.290 437.920 44.890 439.125 ;
        RECT 45.730 437.920 48.110 439.125 ;
        RECT 48.950 437.920 54.550 439.125 ;
        RECT 55.390 437.920 60.990 439.125 ;
        RECT 61.830 437.920 67.430 439.125 ;
        RECT 68.270 437.920 73.870 439.125 ;
        RECT 74.710 437.920 77.090 439.125 ;
        RECT 77.930 437.920 83.530 439.125 ;
        RECT 84.370 437.920 89.970 439.125 ;
        RECT 90.810 437.920 96.410 439.125 ;
        RECT 97.250 437.920 102.850 439.125 ;
        RECT 103.690 437.920 106.070 439.125 ;
        RECT 106.910 437.920 112.510 439.125 ;
        RECT 113.350 437.920 118.950 439.125 ;
        RECT 119.790 437.920 125.390 439.125 ;
        RECT 126.230 437.920 131.830 439.125 ;
        RECT 132.670 437.920 135.050 439.125 ;
        RECT 135.890 437.920 141.490 439.125 ;
        RECT 142.330 437.920 147.930 439.125 ;
        RECT 148.770 437.920 154.370 439.125 ;
        RECT 155.210 437.920 160.810 439.125 ;
        RECT 161.650 437.920 167.250 439.125 ;
        RECT 168.090 437.920 170.470 439.125 ;
        RECT 171.310 437.920 176.910 439.125 ;
        RECT 177.750 437.920 183.350 439.125 ;
        RECT 184.190 437.920 189.790 439.125 ;
        RECT 190.630 437.920 196.230 439.125 ;
        RECT 197.070 437.920 199.450 439.125 ;
        RECT 200.290 437.920 205.890 439.125 ;
        RECT 206.730 437.920 212.330 439.125 ;
        RECT 213.170 437.920 218.770 439.125 ;
        RECT 219.610 437.920 225.210 439.125 ;
        RECT 226.050 437.920 228.430 439.125 ;
        RECT 229.270 437.920 234.870 439.125 ;
        RECT 235.710 437.920 241.310 439.125 ;
        RECT 242.150 437.920 247.750 439.125 ;
        RECT 248.590 437.920 254.190 439.125 ;
        RECT 255.030 437.920 257.410 439.125 ;
        RECT 258.250 437.920 263.850 439.125 ;
        RECT 264.690 437.920 270.290 439.125 ;
        RECT 271.130 437.920 276.730 439.125 ;
        RECT 277.570 437.920 283.170 439.125 ;
        RECT 284.010 437.920 286.390 439.125 ;
        RECT 287.230 437.920 292.830 439.125 ;
        RECT 293.670 437.920 299.270 439.125 ;
        RECT 300.110 437.920 305.710 439.125 ;
        RECT 306.550 437.920 312.150 439.125 ;
        RECT 312.990 437.920 315.370 439.125 ;
        RECT 316.210 437.920 321.810 439.125 ;
        RECT 322.650 437.920 328.250 439.125 ;
        RECT 329.090 437.920 334.690 439.125 ;
        RECT 335.530 437.920 341.130 439.125 ;
        RECT 341.970 437.920 344.350 439.125 ;
        RECT 345.190 437.920 350.790 439.125 ;
        RECT 351.630 437.920 357.230 439.125 ;
        RECT 358.070 437.920 363.670 439.125 ;
        RECT 364.510 437.920 370.110 439.125 ;
        RECT 370.950 437.920 373.330 439.125 ;
        RECT 374.170 437.920 379.770 439.125 ;
        RECT 380.610 437.920 386.210 439.125 ;
        RECT 387.050 437.920 392.650 439.125 ;
        RECT 393.490 437.920 399.090 439.125 ;
        RECT 399.930 437.920 402.310 439.125 ;
        RECT 403.150 437.920 408.750 439.125 ;
        RECT 409.590 437.920 415.190 439.125 ;
        RECT 416.030 437.920 421.630 439.125 ;
        RECT 422.470 437.920 428.070 439.125 ;
        RECT 428.910 437.920 430.460 439.125 ;
        RECT 0.100 4.280 430.460 437.920 ;
        RECT 0.650 3.555 3.030 4.280 ;
        RECT 3.870 3.555 9.470 4.280 ;
        RECT 10.310 3.555 15.910 4.280 ;
        RECT 16.750 3.555 22.350 4.280 ;
        RECT 23.190 3.555 28.790 4.280 ;
        RECT 29.630 3.555 32.010 4.280 ;
        RECT 32.850 3.555 38.450 4.280 ;
        RECT 39.290 3.555 44.890 4.280 ;
        RECT 45.730 3.555 51.330 4.280 ;
        RECT 52.170 3.555 57.770 4.280 ;
        RECT 58.610 3.555 60.990 4.280 ;
        RECT 61.830 3.555 67.430 4.280 ;
        RECT 68.270 3.555 73.870 4.280 ;
        RECT 74.710 3.555 80.310 4.280 ;
        RECT 81.150 3.555 86.750 4.280 ;
        RECT 87.590 3.555 89.970 4.280 ;
        RECT 90.810 3.555 96.410 4.280 ;
        RECT 97.250 3.555 102.850 4.280 ;
        RECT 103.690 3.555 109.290 4.280 ;
        RECT 110.130 3.555 115.730 4.280 ;
        RECT 116.570 3.555 118.950 4.280 ;
        RECT 119.790 3.555 125.390 4.280 ;
        RECT 126.230 3.555 131.830 4.280 ;
        RECT 132.670 3.555 138.270 4.280 ;
        RECT 139.110 3.555 144.710 4.280 ;
        RECT 145.550 3.555 147.930 4.280 ;
        RECT 148.770 3.555 154.370 4.280 ;
        RECT 155.210 3.555 160.810 4.280 ;
        RECT 161.650 3.555 167.250 4.280 ;
        RECT 168.090 3.555 173.690 4.280 ;
        RECT 174.530 3.555 176.910 4.280 ;
        RECT 177.750 3.555 183.350 4.280 ;
        RECT 184.190 3.555 189.790 4.280 ;
        RECT 190.630 3.555 196.230 4.280 ;
        RECT 197.070 3.555 202.670 4.280 ;
        RECT 203.510 3.555 205.890 4.280 ;
        RECT 206.730 3.555 212.330 4.280 ;
        RECT 213.170 3.555 218.770 4.280 ;
        RECT 219.610 3.555 225.210 4.280 ;
        RECT 226.050 3.555 231.650 4.280 ;
        RECT 232.490 3.555 234.870 4.280 ;
        RECT 235.710 3.555 241.310 4.280 ;
        RECT 242.150 3.555 247.750 4.280 ;
        RECT 248.590 3.555 254.190 4.280 ;
        RECT 255.030 3.555 260.630 4.280 ;
        RECT 261.470 3.555 263.850 4.280 ;
        RECT 264.690 3.555 270.290 4.280 ;
        RECT 271.130 3.555 276.730 4.280 ;
        RECT 277.570 3.555 283.170 4.280 ;
        RECT 284.010 3.555 289.610 4.280 ;
        RECT 290.450 3.555 292.830 4.280 ;
        RECT 293.670 3.555 299.270 4.280 ;
        RECT 300.110 3.555 305.710 4.280 ;
        RECT 306.550 3.555 312.150 4.280 ;
        RECT 312.990 3.555 318.590 4.280 ;
        RECT 319.430 3.555 321.810 4.280 ;
        RECT 322.650 3.555 328.250 4.280 ;
        RECT 329.090 3.555 334.690 4.280 ;
        RECT 335.530 3.555 341.130 4.280 ;
        RECT 341.970 3.555 347.570 4.280 ;
        RECT 348.410 3.555 350.790 4.280 ;
        RECT 351.630 3.555 357.230 4.280 ;
        RECT 358.070 3.555 363.670 4.280 ;
        RECT 364.510 3.555 370.110 4.280 ;
        RECT 370.950 3.555 376.550 4.280 ;
        RECT 377.390 3.555 379.770 4.280 ;
        RECT 380.610 3.555 386.210 4.280 ;
        RECT 387.050 3.555 392.650 4.280 ;
        RECT 393.490 3.555 399.090 4.280 ;
        RECT 399.930 3.555 405.530 4.280 ;
        RECT 406.370 3.555 408.750 4.280 ;
        RECT 409.590 3.555 415.190 4.280 ;
        RECT 416.030 3.555 421.630 4.280 ;
        RECT 422.470 3.555 428.070 4.280 ;
        RECT 428.910 3.555 430.460 4.280 ;
      LAYER met3 ;
        RECT 4.400 438.240 427.080 439.105 ;
        RECT 4.000 432.840 428.195 438.240 ;
        RECT 4.400 431.440 427.080 432.840 ;
        RECT 4.000 429.440 428.195 431.440 ;
        RECT 4.400 428.040 428.195 429.440 ;
        RECT 4.000 426.040 428.195 428.040 ;
        RECT 4.000 424.640 427.080 426.040 ;
        RECT 4.000 422.640 428.195 424.640 ;
        RECT 4.400 421.240 428.195 422.640 ;
        RECT 4.000 419.240 428.195 421.240 ;
        RECT 4.000 417.840 427.080 419.240 ;
        RECT 4.000 415.840 428.195 417.840 ;
        RECT 4.400 414.440 428.195 415.840 ;
        RECT 4.000 412.440 428.195 414.440 ;
        RECT 4.000 411.040 427.080 412.440 ;
        RECT 4.000 409.040 428.195 411.040 ;
        RECT 4.400 407.640 427.080 409.040 ;
        RECT 4.000 402.240 428.195 407.640 ;
        RECT 4.400 400.840 427.080 402.240 ;
        RECT 4.000 398.840 428.195 400.840 ;
        RECT 4.400 397.440 428.195 398.840 ;
        RECT 4.000 395.440 428.195 397.440 ;
        RECT 4.000 394.040 427.080 395.440 ;
        RECT 4.000 392.040 428.195 394.040 ;
        RECT 4.400 390.640 428.195 392.040 ;
        RECT 4.000 388.640 428.195 390.640 ;
        RECT 4.000 387.240 427.080 388.640 ;
        RECT 4.000 385.240 428.195 387.240 ;
        RECT 4.400 383.840 428.195 385.240 ;
        RECT 4.000 381.840 428.195 383.840 ;
        RECT 4.000 380.440 427.080 381.840 ;
        RECT 4.000 378.440 428.195 380.440 ;
        RECT 4.400 377.040 427.080 378.440 ;
        RECT 4.000 371.640 428.195 377.040 ;
        RECT 4.400 370.240 427.080 371.640 ;
        RECT 4.000 368.240 428.195 370.240 ;
        RECT 4.400 366.840 428.195 368.240 ;
        RECT 4.000 364.840 428.195 366.840 ;
        RECT 4.000 363.440 427.080 364.840 ;
        RECT 4.000 361.440 428.195 363.440 ;
        RECT 4.400 360.040 428.195 361.440 ;
        RECT 4.000 358.040 428.195 360.040 ;
        RECT 4.000 356.640 427.080 358.040 ;
        RECT 4.000 354.640 428.195 356.640 ;
        RECT 4.400 353.240 428.195 354.640 ;
        RECT 4.000 351.240 428.195 353.240 ;
        RECT 4.000 349.840 427.080 351.240 ;
        RECT 4.000 347.840 428.195 349.840 ;
        RECT 4.400 346.440 427.080 347.840 ;
        RECT 4.000 341.040 428.195 346.440 ;
        RECT 4.400 339.640 427.080 341.040 ;
        RECT 4.000 337.640 428.195 339.640 ;
        RECT 4.400 336.240 428.195 337.640 ;
        RECT 4.000 334.240 428.195 336.240 ;
        RECT 4.000 332.840 427.080 334.240 ;
        RECT 4.000 330.840 428.195 332.840 ;
        RECT 4.400 329.440 428.195 330.840 ;
        RECT 4.000 327.440 428.195 329.440 ;
        RECT 4.000 326.040 427.080 327.440 ;
        RECT 4.000 324.040 428.195 326.040 ;
        RECT 4.400 322.640 428.195 324.040 ;
        RECT 4.000 320.640 428.195 322.640 ;
        RECT 4.000 319.240 427.080 320.640 ;
        RECT 4.000 317.240 428.195 319.240 ;
        RECT 4.400 315.840 427.080 317.240 ;
        RECT 4.000 310.440 428.195 315.840 ;
        RECT 4.400 309.040 427.080 310.440 ;
        RECT 4.000 307.040 428.195 309.040 ;
        RECT 4.400 305.640 428.195 307.040 ;
        RECT 4.000 303.640 428.195 305.640 ;
        RECT 4.000 302.240 427.080 303.640 ;
        RECT 4.000 300.240 428.195 302.240 ;
        RECT 4.400 298.840 428.195 300.240 ;
        RECT 4.000 296.840 428.195 298.840 ;
        RECT 4.000 295.440 427.080 296.840 ;
        RECT 4.000 293.440 428.195 295.440 ;
        RECT 4.400 292.040 428.195 293.440 ;
        RECT 4.000 290.040 428.195 292.040 ;
        RECT 4.000 288.640 427.080 290.040 ;
        RECT 4.000 286.640 428.195 288.640 ;
        RECT 4.400 285.240 427.080 286.640 ;
        RECT 4.000 279.840 428.195 285.240 ;
        RECT 4.400 278.440 427.080 279.840 ;
        RECT 4.000 276.440 428.195 278.440 ;
        RECT 4.400 275.040 428.195 276.440 ;
        RECT 4.000 273.040 428.195 275.040 ;
        RECT 4.000 271.640 427.080 273.040 ;
        RECT 4.000 269.640 428.195 271.640 ;
        RECT 4.400 268.240 428.195 269.640 ;
        RECT 4.000 266.240 428.195 268.240 ;
        RECT 4.000 264.840 427.080 266.240 ;
        RECT 4.000 262.840 428.195 264.840 ;
        RECT 4.400 261.440 428.195 262.840 ;
        RECT 4.000 259.440 428.195 261.440 ;
        RECT 4.000 258.040 427.080 259.440 ;
        RECT 4.000 256.040 428.195 258.040 ;
        RECT 4.400 254.640 427.080 256.040 ;
        RECT 4.000 249.240 428.195 254.640 ;
        RECT 4.400 247.840 427.080 249.240 ;
        RECT 4.000 245.840 428.195 247.840 ;
        RECT 4.400 244.440 428.195 245.840 ;
        RECT 4.000 242.440 428.195 244.440 ;
        RECT 4.000 241.040 427.080 242.440 ;
        RECT 4.000 239.040 428.195 241.040 ;
        RECT 4.400 237.640 428.195 239.040 ;
        RECT 4.000 235.640 428.195 237.640 ;
        RECT 4.000 234.240 427.080 235.640 ;
        RECT 4.000 232.240 428.195 234.240 ;
        RECT 4.400 230.840 428.195 232.240 ;
        RECT 4.000 228.840 428.195 230.840 ;
        RECT 4.000 227.440 427.080 228.840 ;
        RECT 4.000 225.440 428.195 227.440 ;
        RECT 4.400 224.040 427.080 225.440 ;
        RECT 4.000 218.640 428.195 224.040 ;
        RECT 4.400 217.240 427.080 218.640 ;
        RECT 4.000 215.240 428.195 217.240 ;
        RECT 4.400 213.840 428.195 215.240 ;
        RECT 4.000 211.840 428.195 213.840 ;
        RECT 4.000 210.440 427.080 211.840 ;
        RECT 4.000 208.440 428.195 210.440 ;
        RECT 4.400 207.040 428.195 208.440 ;
        RECT 4.000 205.040 428.195 207.040 ;
        RECT 4.000 203.640 427.080 205.040 ;
        RECT 4.000 201.640 428.195 203.640 ;
        RECT 4.400 200.240 428.195 201.640 ;
        RECT 4.000 198.240 428.195 200.240 ;
        RECT 4.000 196.840 427.080 198.240 ;
        RECT 4.000 194.840 428.195 196.840 ;
        RECT 4.400 193.440 427.080 194.840 ;
        RECT 4.000 188.040 428.195 193.440 ;
        RECT 4.400 186.640 427.080 188.040 ;
        RECT 4.000 184.640 428.195 186.640 ;
        RECT 4.400 183.240 428.195 184.640 ;
        RECT 4.000 181.240 428.195 183.240 ;
        RECT 4.000 179.840 427.080 181.240 ;
        RECT 4.000 177.840 428.195 179.840 ;
        RECT 4.400 176.440 428.195 177.840 ;
        RECT 4.000 174.440 428.195 176.440 ;
        RECT 4.000 173.040 427.080 174.440 ;
        RECT 4.000 171.040 428.195 173.040 ;
        RECT 4.400 169.640 428.195 171.040 ;
        RECT 4.000 167.640 428.195 169.640 ;
        RECT 4.000 166.240 427.080 167.640 ;
        RECT 4.000 164.240 428.195 166.240 ;
        RECT 4.400 162.840 427.080 164.240 ;
        RECT 4.000 157.440 428.195 162.840 ;
        RECT 4.400 156.040 427.080 157.440 ;
        RECT 4.000 154.040 428.195 156.040 ;
        RECT 4.400 152.640 428.195 154.040 ;
        RECT 4.000 150.640 428.195 152.640 ;
        RECT 4.000 149.240 427.080 150.640 ;
        RECT 4.000 147.240 428.195 149.240 ;
        RECT 4.400 145.840 428.195 147.240 ;
        RECT 4.000 143.840 428.195 145.840 ;
        RECT 4.000 142.440 427.080 143.840 ;
        RECT 4.000 140.440 428.195 142.440 ;
        RECT 4.400 139.040 428.195 140.440 ;
        RECT 4.000 137.040 428.195 139.040 ;
        RECT 4.000 135.640 427.080 137.040 ;
        RECT 4.000 133.640 428.195 135.640 ;
        RECT 4.400 132.240 428.195 133.640 ;
        RECT 4.000 130.240 428.195 132.240 ;
        RECT 4.000 128.840 427.080 130.240 ;
        RECT 4.000 126.840 428.195 128.840 ;
        RECT 4.400 125.440 427.080 126.840 ;
        RECT 4.000 123.440 428.195 125.440 ;
        RECT 4.400 122.040 428.195 123.440 ;
        RECT 4.000 120.040 428.195 122.040 ;
        RECT 4.000 118.640 427.080 120.040 ;
        RECT 4.000 116.640 428.195 118.640 ;
        RECT 4.400 115.240 428.195 116.640 ;
        RECT 4.000 113.240 428.195 115.240 ;
        RECT 4.000 111.840 427.080 113.240 ;
        RECT 4.000 109.840 428.195 111.840 ;
        RECT 4.400 108.440 428.195 109.840 ;
        RECT 4.000 106.440 428.195 108.440 ;
        RECT 4.000 105.040 427.080 106.440 ;
        RECT 4.000 103.040 428.195 105.040 ;
        RECT 4.400 101.640 428.195 103.040 ;
        RECT 4.000 99.640 428.195 101.640 ;
        RECT 4.000 98.240 427.080 99.640 ;
        RECT 4.000 96.240 428.195 98.240 ;
        RECT 4.400 94.840 427.080 96.240 ;
        RECT 4.000 92.840 428.195 94.840 ;
        RECT 4.400 91.440 428.195 92.840 ;
        RECT 4.000 89.440 428.195 91.440 ;
        RECT 4.000 88.040 427.080 89.440 ;
        RECT 4.000 86.040 428.195 88.040 ;
        RECT 4.400 84.640 428.195 86.040 ;
        RECT 4.000 82.640 428.195 84.640 ;
        RECT 4.000 81.240 427.080 82.640 ;
        RECT 4.000 79.240 428.195 81.240 ;
        RECT 4.400 77.840 428.195 79.240 ;
        RECT 4.000 75.840 428.195 77.840 ;
        RECT 4.000 74.440 427.080 75.840 ;
        RECT 4.000 72.440 428.195 74.440 ;
        RECT 4.400 71.040 428.195 72.440 ;
        RECT 4.000 69.040 428.195 71.040 ;
        RECT 4.000 67.640 427.080 69.040 ;
        RECT 4.000 65.640 428.195 67.640 ;
        RECT 4.400 64.240 427.080 65.640 ;
        RECT 4.000 62.240 428.195 64.240 ;
        RECT 4.400 60.840 428.195 62.240 ;
        RECT 4.000 58.840 428.195 60.840 ;
        RECT 4.000 57.440 427.080 58.840 ;
        RECT 4.000 55.440 428.195 57.440 ;
        RECT 4.400 54.040 428.195 55.440 ;
        RECT 4.000 52.040 428.195 54.040 ;
        RECT 4.000 50.640 427.080 52.040 ;
        RECT 4.000 48.640 428.195 50.640 ;
        RECT 4.400 47.240 428.195 48.640 ;
        RECT 4.000 45.240 428.195 47.240 ;
        RECT 4.000 43.840 427.080 45.240 ;
        RECT 4.000 41.840 428.195 43.840 ;
        RECT 4.400 40.440 428.195 41.840 ;
        RECT 4.000 38.440 428.195 40.440 ;
        RECT 4.000 37.040 427.080 38.440 ;
        RECT 4.000 35.040 428.195 37.040 ;
        RECT 4.400 33.640 427.080 35.040 ;
        RECT 4.000 31.640 428.195 33.640 ;
        RECT 4.400 30.240 428.195 31.640 ;
        RECT 4.000 28.240 428.195 30.240 ;
        RECT 4.000 26.840 427.080 28.240 ;
        RECT 4.000 24.840 428.195 26.840 ;
        RECT 4.400 23.440 428.195 24.840 ;
        RECT 4.000 21.440 428.195 23.440 ;
        RECT 4.000 20.040 427.080 21.440 ;
        RECT 4.000 18.040 428.195 20.040 ;
        RECT 4.400 16.640 428.195 18.040 ;
        RECT 4.000 14.640 428.195 16.640 ;
        RECT 4.000 13.240 427.080 14.640 ;
        RECT 4.000 11.240 428.195 13.240 ;
        RECT 4.400 9.840 428.195 11.240 ;
        RECT 4.000 7.840 428.195 9.840 ;
        RECT 4.000 6.440 427.080 7.840 ;
        RECT 4.000 4.440 428.195 6.440 ;
        RECT 4.400 3.575 427.080 4.440 ;
      LAYER met4 ;
        RECT 33.415 430.400 419.225 431.625 ;
        RECT 33.415 10.240 174.240 430.400 ;
        RECT 176.640 10.240 177.540 430.400 ;
        RECT 179.940 10.240 327.840 430.400 ;
        RECT 330.240 10.240 331.140 430.400 ;
        RECT 333.540 10.240 419.225 430.400 ;
        RECT 33.415 9.695 419.225 10.240 ;
      LAYER met5 ;
        RECT 113.740 119.900 181.580 121.500 ;
  END
END password_cracker
END LIBRARY

