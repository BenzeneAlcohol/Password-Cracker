module password_cracker (clk,
    cracked,
    done,
    init,
    reset,
    VPWR,
    VGND,
    hash,
    password_count);
 input clk;
 output cracked;
 output done;
 input init;
 input reset;
 input VPWR;
 input VGND;
 input [255:0] hash;
 output [31:0] password_count;

 wire Hash_Digest;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire net261;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net262;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net263;
 wire net291;
 wire clknet_leaf_0_clk;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire \sha256cu.K[0] ;
 wire \sha256cu.K[10] ;
 wire \sha256cu.K[11] ;
 wire \sha256cu.K[12] ;
 wire \sha256cu.K[13] ;
 wire \sha256cu.K[14] ;
 wire \sha256cu.K[15] ;
 wire \sha256cu.K[16] ;
 wire \sha256cu.K[17] ;
 wire \sha256cu.K[18] ;
 wire \sha256cu.K[19] ;
 wire \sha256cu.K[1] ;
 wire \sha256cu.K[20] ;
 wire \sha256cu.K[21] ;
 wire \sha256cu.K[22] ;
 wire \sha256cu.K[23] ;
 wire \sha256cu.K[24] ;
 wire \sha256cu.K[25] ;
 wire \sha256cu.K[26] ;
 wire \sha256cu.K[27] ;
 wire \sha256cu.K[28] ;
 wire \sha256cu.K[29] ;
 wire \sha256cu.K[2] ;
 wire \sha256cu.K[30] ;
 wire \sha256cu.K[31] ;
 wire \sha256cu.K[3] ;
 wire \sha256cu.K[4] ;
 wire \sha256cu.K[5] ;
 wire \sha256cu.K[6] ;
 wire \sha256cu.K[7] ;
 wire \sha256cu.K[8] ;
 wire \sha256cu.K[9] ;
 wire \sha256cu.byte_rdy ;
 wire \sha256cu.byte_stop ;
 wire \sha256cu.counter_iteration[0] ;
 wire \sha256cu.counter_iteration[1] ;
 wire \sha256cu.counter_iteration[2] ;
 wire \sha256cu.counter_iteration[3] ;
 wire \sha256cu.counter_iteration[4] ;
 wire \sha256cu.counter_iteration[5] ;
 wire \sha256cu.counter_iteration[6] ;
 wire \sha256cu.data_in_padd[0] ;
 wire \sha256cu.data_in_padd[10] ;
 wire \sha256cu.data_in_padd[11] ;
 wire \sha256cu.data_in_padd[12] ;
 wire \sha256cu.data_in_padd[13] ;
 wire \sha256cu.data_in_padd[14] ;
 wire \sha256cu.data_in_padd[15] ;
 wire \sha256cu.data_in_padd[16] ;
 wire \sha256cu.data_in_padd[17] ;
 wire \sha256cu.data_in_padd[18] ;
 wire \sha256cu.data_in_padd[19] ;
 wire \sha256cu.data_in_padd[1] ;
 wire \sha256cu.data_in_padd[20] ;
 wire \sha256cu.data_in_padd[21] ;
 wire \sha256cu.data_in_padd[22] ;
 wire \sha256cu.data_in_padd[23] ;
 wire \sha256cu.data_in_padd[24] ;
 wire \sha256cu.data_in_padd[25] ;
 wire \sha256cu.data_in_padd[26] ;
 wire \sha256cu.data_in_padd[27] ;
 wire \sha256cu.data_in_padd[28] ;
 wire \sha256cu.data_in_padd[29] ;
 wire \sha256cu.data_in_padd[2] ;
 wire \sha256cu.data_in_padd[30] ;
 wire \sha256cu.data_in_padd[31] ;
 wire \sha256cu.data_in_padd[3] ;
 wire \sha256cu.data_in_padd[4] ;
 wire \sha256cu.data_in_padd[5] ;
 wire \sha256cu.data_in_padd[6] ;
 wire \sha256cu.data_in_padd[7] ;
 wire \sha256cu.data_in_padd[8] ;
 wire \sha256cu.data_in_padd[9] ;
 wire \sha256cu.flag_0_15 ;
 wire \sha256cu.hashing_done ;
 wire \sha256cu.iter_processing.padding_done ;
 wire \sha256cu.iter_processing.rst ;
 wire \sha256cu.iter_processing.temp_case ;
 wire \sha256cu.iter_processing.temp_if ;
 wire \sha256cu.iter_processing.w[0] ;
 wire \sha256cu.iter_processing.w[10] ;
 wire \sha256cu.iter_processing.w[11] ;
 wire \sha256cu.iter_processing.w[12] ;
 wire \sha256cu.iter_processing.w[13] ;
 wire \sha256cu.iter_processing.w[14] ;
 wire \sha256cu.iter_processing.w[15] ;
 wire \sha256cu.iter_processing.w[16] ;
 wire \sha256cu.iter_processing.w[17] ;
 wire \sha256cu.iter_processing.w[18] ;
 wire \sha256cu.iter_processing.w[19] ;
 wire \sha256cu.iter_processing.w[1] ;
 wire \sha256cu.iter_processing.w[20] ;
 wire \sha256cu.iter_processing.w[21] ;
 wire \sha256cu.iter_processing.w[22] ;
 wire \sha256cu.iter_processing.w[23] ;
 wire \sha256cu.iter_processing.w[24] ;
 wire \sha256cu.iter_processing.w[25] ;
 wire \sha256cu.iter_processing.w[26] ;
 wire \sha256cu.iter_processing.w[27] ;
 wire \sha256cu.iter_processing.w[28] ;
 wire \sha256cu.iter_processing.w[29] ;
 wire \sha256cu.iter_processing.w[2] ;
 wire \sha256cu.iter_processing.w[30] ;
 wire \sha256cu.iter_processing.w[31] ;
 wire \sha256cu.iter_processing.w[3] ;
 wire \sha256cu.iter_processing.w[4] ;
 wire \sha256cu.iter_processing.w[5] ;
 wire \sha256cu.iter_processing.w[6] ;
 wire \sha256cu.iter_processing.w[7] ;
 wire \sha256cu.iter_processing.w[8] ;
 wire \sha256cu.iter_processing.w[9] ;
 wire \sha256cu.m_out_digest.H7[0] ;
 wire \sha256cu.m_out_digest.a_in[0] ;
 wire \sha256cu.m_out_digest.a_in[10] ;
 wire \sha256cu.m_out_digest.a_in[11] ;
 wire \sha256cu.m_out_digest.a_in[12] ;
 wire \sha256cu.m_out_digest.a_in[13] ;
 wire \sha256cu.m_out_digest.a_in[14] ;
 wire \sha256cu.m_out_digest.a_in[15] ;
 wire \sha256cu.m_out_digest.a_in[16] ;
 wire \sha256cu.m_out_digest.a_in[17] ;
 wire \sha256cu.m_out_digest.a_in[18] ;
 wire \sha256cu.m_out_digest.a_in[19] ;
 wire \sha256cu.m_out_digest.a_in[1] ;
 wire \sha256cu.m_out_digest.a_in[20] ;
 wire \sha256cu.m_out_digest.a_in[21] ;
 wire \sha256cu.m_out_digest.a_in[22] ;
 wire \sha256cu.m_out_digest.a_in[23] ;
 wire \sha256cu.m_out_digest.a_in[24] ;
 wire \sha256cu.m_out_digest.a_in[25] ;
 wire \sha256cu.m_out_digest.a_in[26] ;
 wire \sha256cu.m_out_digest.a_in[27] ;
 wire \sha256cu.m_out_digest.a_in[28] ;
 wire \sha256cu.m_out_digest.a_in[29] ;
 wire \sha256cu.m_out_digest.a_in[2] ;
 wire \sha256cu.m_out_digest.a_in[30] ;
 wire \sha256cu.m_out_digest.a_in[31] ;
 wire \sha256cu.m_out_digest.a_in[3] ;
 wire \sha256cu.m_out_digest.a_in[4] ;
 wire \sha256cu.m_out_digest.a_in[5] ;
 wire \sha256cu.m_out_digest.a_in[6] ;
 wire \sha256cu.m_out_digest.a_in[7] ;
 wire \sha256cu.m_out_digest.a_in[8] ;
 wire \sha256cu.m_out_digest.a_in[9] ;
 wire \sha256cu.m_out_digest.b_in[0] ;
 wire \sha256cu.m_out_digest.b_in[10] ;
 wire \sha256cu.m_out_digest.b_in[11] ;
 wire \sha256cu.m_out_digest.b_in[12] ;
 wire \sha256cu.m_out_digest.b_in[13] ;
 wire \sha256cu.m_out_digest.b_in[14] ;
 wire \sha256cu.m_out_digest.b_in[15] ;
 wire \sha256cu.m_out_digest.b_in[16] ;
 wire \sha256cu.m_out_digest.b_in[17] ;
 wire \sha256cu.m_out_digest.b_in[18] ;
 wire \sha256cu.m_out_digest.b_in[19] ;
 wire \sha256cu.m_out_digest.b_in[1] ;
 wire \sha256cu.m_out_digest.b_in[20] ;
 wire \sha256cu.m_out_digest.b_in[21] ;
 wire \sha256cu.m_out_digest.b_in[22] ;
 wire \sha256cu.m_out_digest.b_in[23] ;
 wire \sha256cu.m_out_digest.b_in[24] ;
 wire \sha256cu.m_out_digest.b_in[25] ;
 wire \sha256cu.m_out_digest.b_in[26] ;
 wire \sha256cu.m_out_digest.b_in[27] ;
 wire \sha256cu.m_out_digest.b_in[28] ;
 wire \sha256cu.m_out_digest.b_in[29] ;
 wire \sha256cu.m_out_digest.b_in[2] ;
 wire \sha256cu.m_out_digest.b_in[30] ;
 wire \sha256cu.m_out_digest.b_in[31] ;
 wire \sha256cu.m_out_digest.b_in[3] ;
 wire \sha256cu.m_out_digest.b_in[4] ;
 wire \sha256cu.m_out_digest.b_in[5] ;
 wire \sha256cu.m_out_digest.b_in[6] ;
 wire \sha256cu.m_out_digest.b_in[7] ;
 wire \sha256cu.m_out_digest.b_in[8] ;
 wire \sha256cu.m_out_digest.b_in[9] ;
 wire \sha256cu.m_out_digest.c_in[0] ;
 wire \sha256cu.m_out_digest.c_in[10] ;
 wire \sha256cu.m_out_digest.c_in[11] ;
 wire \sha256cu.m_out_digest.c_in[12] ;
 wire \sha256cu.m_out_digest.c_in[13] ;
 wire \sha256cu.m_out_digest.c_in[14] ;
 wire \sha256cu.m_out_digest.c_in[15] ;
 wire \sha256cu.m_out_digest.c_in[16] ;
 wire \sha256cu.m_out_digest.c_in[17] ;
 wire \sha256cu.m_out_digest.c_in[18] ;
 wire \sha256cu.m_out_digest.c_in[19] ;
 wire \sha256cu.m_out_digest.c_in[1] ;
 wire \sha256cu.m_out_digest.c_in[20] ;
 wire \sha256cu.m_out_digest.c_in[21] ;
 wire \sha256cu.m_out_digest.c_in[22] ;
 wire \sha256cu.m_out_digest.c_in[23] ;
 wire \sha256cu.m_out_digest.c_in[24] ;
 wire \sha256cu.m_out_digest.c_in[25] ;
 wire \sha256cu.m_out_digest.c_in[26] ;
 wire \sha256cu.m_out_digest.c_in[27] ;
 wire \sha256cu.m_out_digest.c_in[28] ;
 wire \sha256cu.m_out_digest.c_in[29] ;
 wire \sha256cu.m_out_digest.c_in[2] ;
 wire \sha256cu.m_out_digest.c_in[30] ;
 wire \sha256cu.m_out_digest.c_in[31] ;
 wire \sha256cu.m_out_digest.c_in[3] ;
 wire \sha256cu.m_out_digest.c_in[4] ;
 wire \sha256cu.m_out_digest.c_in[5] ;
 wire \sha256cu.m_out_digest.c_in[6] ;
 wire \sha256cu.m_out_digest.c_in[7] ;
 wire \sha256cu.m_out_digest.c_in[8] ;
 wire \sha256cu.m_out_digest.c_in[9] ;
 wire \sha256cu.m_out_digest.d_in[0] ;
 wire \sha256cu.m_out_digest.d_in[10] ;
 wire \sha256cu.m_out_digest.d_in[11] ;
 wire \sha256cu.m_out_digest.d_in[12] ;
 wire \sha256cu.m_out_digest.d_in[13] ;
 wire \sha256cu.m_out_digest.d_in[14] ;
 wire \sha256cu.m_out_digest.d_in[15] ;
 wire \sha256cu.m_out_digest.d_in[16] ;
 wire \sha256cu.m_out_digest.d_in[17] ;
 wire \sha256cu.m_out_digest.d_in[18] ;
 wire \sha256cu.m_out_digest.d_in[19] ;
 wire \sha256cu.m_out_digest.d_in[1] ;
 wire \sha256cu.m_out_digest.d_in[20] ;
 wire \sha256cu.m_out_digest.d_in[21] ;
 wire \sha256cu.m_out_digest.d_in[22] ;
 wire \sha256cu.m_out_digest.d_in[23] ;
 wire \sha256cu.m_out_digest.d_in[24] ;
 wire \sha256cu.m_out_digest.d_in[25] ;
 wire \sha256cu.m_out_digest.d_in[26] ;
 wire \sha256cu.m_out_digest.d_in[27] ;
 wire \sha256cu.m_out_digest.d_in[28] ;
 wire \sha256cu.m_out_digest.d_in[29] ;
 wire \sha256cu.m_out_digest.d_in[2] ;
 wire \sha256cu.m_out_digest.d_in[30] ;
 wire \sha256cu.m_out_digest.d_in[31] ;
 wire \sha256cu.m_out_digest.d_in[3] ;
 wire \sha256cu.m_out_digest.d_in[4] ;
 wire \sha256cu.m_out_digest.d_in[5] ;
 wire \sha256cu.m_out_digest.d_in[6] ;
 wire \sha256cu.m_out_digest.d_in[7] ;
 wire \sha256cu.m_out_digest.d_in[8] ;
 wire \sha256cu.m_out_digest.d_in[9] ;
 wire \sha256cu.m_out_digest.e_in[0] ;
 wire \sha256cu.m_out_digest.e_in[10] ;
 wire \sha256cu.m_out_digest.e_in[11] ;
 wire \sha256cu.m_out_digest.e_in[12] ;
 wire \sha256cu.m_out_digest.e_in[13] ;
 wire \sha256cu.m_out_digest.e_in[14] ;
 wire \sha256cu.m_out_digest.e_in[15] ;
 wire \sha256cu.m_out_digest.e_in[16] ;
 wire \sha256cu.m_out_digest.e_in[17] ;
 wire \sha256cu.m_out_digest.e_in[18] ;
 wire \sha256cu.m_out_digest.e_in[19] ;
 wire \sha256cu.m_out_digest.e_in[1] ;
 wire \sha256cu.m_out_digest.e_in[20] ;
 wire \sha256cu.m_out_digest.e_in[21] ;
 wire \sha256cu.m_out_digest.e_in[22] ;
 wire \sha256cu.m_out_digest.e_in[23] ;
 wire \sha256cu.m_out_digest.e_in[24] ;
 wire \sha256cu.m_out_digest.e_in[25] ;
 wire \sha256cu.m_out_digest.e_in[26] ;
 wire \sha256cu.m_out_digest.e_in[27] ;
 wire \sha256cu.m_out_digest.e_in[28] ;
 wire \sha256cu.m_out_digest.e_in[29] ;
 wire \sha256cu.m_out_digest.e_in[2] ;
 wire \sha256cu.m_out_digest.e_in[30] ;
 wire \sha256cu.m_out_digest.e_in[31] ;
 wire \sha256cu.m_out_digest.e_in[3] ;
 wire \sha256cu.m_out_digest.e_in[4] ;
 wire \sha256cu.m_out_digest.e_in[5] ;
 wire \sha256cu.m_out_digest.e_in[6] ;
 wire \sha256cu.m_out_digest.e_in[7] ;
 wire \sha256cu.m_out_digest.e_in[8] ;
 wire \sha256cu.m_out_digest.e_in[9] ;
 wire \sha256cu.m_out_digest.f_in[0] ;
 wire \sha256cu.m_out_digest.f_in[10] ;
 wire \sha256cu.m_out_digest.f_in[11] ;
 wire \sha256cu.m_out_digest.f_in[12] ;
 wire \sha256cu.m_out_digest.f_in[13] ;
 wire \sha256cu.m_out_digest.f_in[14] ;
 wire \sha256cu.m_out_digest.f_in[15] ;
 wire \sha256cu.m_out_digest.f_in[16] ;
 wire \sha256cu.m_out_digest.f_in[17] ;
 wire \sha256cu.m_out_digest.f_in[18] ;
 wire \sha256cu.m_out_digest.f_in[19] ;
 wire \sha256cu.m_out_digest.f_in[1] ;
 wire \sha256cu.m_out_digest.f_in[20] ;
 wire \sha256cu.m_out_digest.f_in[21] ;
 wire \sha256cu.m_out_digest.f_in[22] ;
 wire \sha256cu.m_out_digest.f_in[23] ;
 wire \sha256cu.m_out_digest.f_in[24] ;
 wire \sha256cu.m_out_digest.f_in[25] ;
 wire \sha256cu.m_out_digest.f_in[26] ;
 wire \sha256cu.m_out_digest.f_in[27] ;
 wire \sha256cu.m_out_digest.f_in[28] ;
 wire \sha256cu.m_out_digest.f_in[29] ;
 wire \sha256cu.m_out_digest.f_in[2] ;
 wire \sha256cu.m_out_digest.f_in[30] ;
 wire \sha256cu.m_out_digest.f_in[31] ;
 wire \sha256cu.m_out_digest.f_in[3] ;
 wire \sha256cu.m_out_digest.f_in[4] ;
 wire \sha256cu.m_out_digest.f_in[5] ;
 wire \sha256cu.m_out_digest.f_in[6] ;
 wire \sha256cu.m_out_digest.f_in[7] ;
 wire \sha256cu.m_out_digest.f_in[8] ;
 wire \sha256cu.m_out_digest.f_in[9] ;
 wire \sha256cu.m_out_digest.g_in[0] ;
 wire \sha256cu.m_out_digest.g_in[10] ;
 wire \sha256cu.m_out_digest.g_in[11] ;
 wire \sha256cu.m_out_digest.g_in[12] ;
 wire \sha256cu.m_out_digest.g_in[13] ;
 wire \sha256cu.m_out_digest.g_in[14] ;
 wire \sha256cu.m_out_digest.g_in[15] ;
 wire \sha256cu.m_out_digest.g_in[16] ;
 wire \sha256cu.m_out_digest.g_in[17] ;
 wire \sha256cu.m_out_digest.g_in[18] ;
 wire \sha256cu.m_out_digest.g_in[19] ;
 wire \sha256cu.m_out_digest.g_in[1] ;
 wire \sha256cu.m_out_digest.g_in[20] ;
 wire \sha256cu.m_out_digest.g_in[21] ;
 wire \sha256cu.m_out_digest.g_in[22] ;
 wire \sha256cu.m_out_digest.g_in[23] ;
 wire \sha256cu.m_out_digest.g_in[24] ;
 wire \sha256cu.m_out_digest.g_in[25] ;
 wire \sha256cu.m_out_digest.g_in[26] ;
 wire \sha256cu.m_out_digest.g_in[27] ;
 wire \sha256cu.m_out_digest.g_in[28] ;
 wire \sha256cu.m_out_digest.g_in[29] ;
 wire \sha256cu.m_out_digest.g_in[2] ;
 wire \sha256cu.m_out_digest.g_in[30] ;
 wire \sha256cu.m_out_digest.g_in[31] ;
 wire \sha256cu.m_out_digest.g_in[3] ;
 wire \sha256cu.m_out_digest.g_in[4] ;
 wire \sha256cu.m_out_digest.g_in[5] ;
 wire \sha256cu.m_out_digest.g_in[6] ;
 wire \sha256cu.m_out_digest.g_in[7] ;
 wire \sha256cu.m_out_digest.g_in[8] ;
 wire \sha256cu.m_out_digest.g_in[9] ;
 wire \sha256cu.m_out_digest.h_in[0] ;
 wire \sha256cu.m_out_digest.h_in[10] ;
 wire \sha256cu.m_out_digest.h_in[11] ;
 wire \sha256cu.m_out_digest.h_in[12] ;
 wire \sha256cu.m_out_digest.h_in[13] ;
 wire \sha256cu.m_out_digest.h_in[14] ;
 wire \sha256cu.m_out_digest.h_in[15] ;
 wire \sha256cu.m_out_digest.h_in[16] ;
 wire \sha256cu.m_out_digest.h_in[17] ;
 wire \sha256cu.m_out_digest.h_in[18] ;
 wire \sha256cu.m_out_digest.h_in[19] ;
 wire \sha256cu.m_out_digest.h_in[1] ;
 wire \sha256cu.m_out_digest.h_in[20] ;
 wire \sha256cu.m_out_digest.h_in[21] ;
 wire \sha256cu.m_out_digest.h_in[22] ;
 wire \sha256cu.m_out_digest.h_in[23] ;
 wire \sha256cu.m_out_digest.h_in[24] ;
 wire \sha256cu.m_out_digest.h_in[25] ;
 wire \sha256cu.m_out_digest.h_in[26] ;
 wire \sha256cu.m_out_digest.h_in[27] ;
 wire \sha256cu.m_out_digest.h_in[28] ;
 wire \sha256cu.m_out_digest.h_in[29] ;
 wire \sha256cu.m_out_digest.h_in[2] ;
 wire \sha256cu.m_out_digest.h_in[30] ;
 wire \sha256cu.m_out_digest.h_in[31] ;
 wire \sha256cu.m_out_digest.h_in[3] ;
 wire \sha256cu.m_out_digest.h_in[4] ;
 wire \sha256cu.m_out_digest.h_in[5] ;
 wire \sha256cu.m_out_digest.h_in[6] ;
 wire \sha256cu.m_out_digest.h_in[7] ;
 wire \sha256cu.m_out_digest.h_in[8] ;
 wire \sha256cu.m_out_digest.h_in[9] ;
 wire \sha256cu.m_out_digest.temp_delay ;
 wire \sha256cu.m_pad_pars.add_512_block[0] ;
 wire \sha256cu.m_pad_pars.add_512_block[1] ;
 wire \sha256cu.m_pad_pars.add_512_block[2] ;
 wire \sha256cu.m_pad_pars.add_512_block[3] ;
 wire \sha256cu.m_pad_pars.add_512_block[4] ;
 wire \sha256cu.m_pad_pars.add_512_block[5] ;
 wire \sha256cu.m_pad_pars.add_512_block[6] ;
 wire \sha256cu.m_pad_pars.add_out0[2] ;
 wire \sha256cu.m_pad_pars.add_out0[3] ;
 wire \sha256cu.m_pad_pars.add_out0[4] ;
 wire \sha256cu.m_pad_pars.add_out0[5] ;
 wire \sha256cu.m_pad_pars.add_out0[6] ;
 wire \sha256cu.m_pad_pars.add_out1[2] ;
 wire \sha256cu.m_pad_pars.add_out1[3] ;
 wire \sha256cu.m_pad_pars.add_out1[4] ;
 wire \sha256cu.m_pad_pars.add_out1[5] ;
 wire \sha256cu.m_pad_pars.add_out2[2] ;
 wire \sha256cu.m_pad_pars.add_out2[3] ;
 wire \sha256cu.m_pad_pars.add_out2[4] ;
 wire \sha256cu.m_pad_pars.add_out2[5] ;
 wire \sha256cu.m_pad_pars.add_out3[2] ;
 wire \sha256cu.m_pad_pars.add_out3[3] ;
 wire \sha256cu.m_pad_pars.add_out3[4] ;
 wire \sha256cu.m_pad_pars.add_out3[5] ;
 wire \sha256cu.m_pad_pars.add_out3[6] ;
 wire \sha256cu.m_pad_pars.block_512[0][0] ;
 wire \sha256cu.m_pad_pars.block_512[0][1] ;
 wire \sha256cu.m_pad_pars.block_512[0][2] ;
 wire \sha256cu.m_pad_pars.block_512[0][3] ;
 wire \sha256cu.m_pad_pars.block_512[0][4] ;
 wire \sha256cu.m_pad_pars.block_512[0][5] ;
 wire \sha256cu.m_pad_pars.block_512[0][6] ;
 wire \sha256cu.m_pad_pars.block_512[0][7] ;
 wire \sha256cu.m_pad_pars.block_512[10][0] ;
 wire \sha256cu.m_pad_pars.block_512[10][1] ;
 wire \sha256cu.m_pad_pars.block_512[10][2] ;
 wire \sha256cu.m_pad_pars.block_512[10][3] ;
 wire \sha256cu.m_pad_pars.block_512[10][4] ;
 wire \sha256cu.m_pad_pars.block_512[10][5] ;
 wire \sha256cu.m_pad_pars.block_512[10][6] ;
 wire \sha256cu.m_pad_pars.block_512[10][7] ;
 wire \sha256cu.m_pad_pars.block_512[11][0] ;
 wire \sha256cu.m_pad_pars.block_512[11][1] ;
 wire \sha256cu.m_pad_pars.block_512[11][2] ;
 wire \sha256cu.m_pad_pars.block_512[11][3] ;
 wire \sha256cu.m_pad_pars.block_512[11][4] ;
 wire \sha256cu.m_pad_pars.block_512[11][5] ;
 wire \sha256cu.m_pad_pars.block_512[11][6] ;
 wire \sha256cu.m_pad_pars.block_512[11][7] ;
 wire \sha256cu.m_pad_pars.block_512[12][0] ;
 wire \sha256cu.m_pad_pars.block_512[12][1] ;
 wire \sha256cu.m_pad_pars.block_512[12][2] ;
 wire \sha256cu.m_pad_pars.block_512[12][3] ;
 wire \sha256cu.m_pad_pars.block_512[12][4] ;
 wire \sha256cu.m_pad_pars.block_512[12][5] ;
 wire \sha256cu.m_pad_pars.block_512[12][6] ;
 wire \sha256cu.m_pad_pars.block_512[12][7] ;
 wire \sha256cu.m_pad_pars.block_512[13][0] ;
 wire \sha256cu.m_pad_pars.block_512[13][1] ;
 wire \sha256cu.m_pad_pars.block_512[13][2] ;
 wire \sha256cu.m_pad_pars.block_512[13][3] ;
 wire \sha256cu.m_pad_pars.block_512[13][4] ;
 wire \sha256cu.m_pad_pars.block_512[13][5] ;
 wire \sha256cu.m_pad_pars.block_512[13][6] ;
 wire \sha256cu.m_pad_pars.block_512[13][7] ;
 wire \sha256cu.m_pad_pars.block_512[14][0] ;
 wire \sha256cu.m_pad_pars.block_512[14][1] ;
 wire \sha256cu.m_pad_pars.block_512[14][2] ;
 wire \sha256cu.m_pad_pars.block_512[14][3] ;
 wire \sha256cu.m_pad_pars.block_512[14][4] ;
 wire \sha256cu.m_pad_pars.block_512[14][5] ;
 wire \sha256cu.m_pad_pars.block_512[14][6] ;
 wire \sha256cu.m_pad_pars.block_512[14][7] ;
 wire \sha256cu.m_pad_pars.block_512[15][0] ;
 wire \sha256cu.m_pad_pars.block_512[15][1] ;
 wire \sha256cu.m_pad_pars.block_512[15][2] ;
 wire \sha256cu.m_pad_pars.block_512[15][3] ;
 wire \sha256cu.m_pad_pars.block_512[15][4] ;
 wire \sha256cu.m_pad_pars.block_512[15][5] ;
 wire \sha256cu.m_pad_pars.block_512[15][6] ;
 wire \sha256cu.m_pad_pars.block_512[15][7] ;
 wire \sha256cu.m_pad_pars.block_512[16][0] ;
 wire \sha256cu.m_pad_pars.block_512[16][1] ;
 wire \sha256cu.m_pad_pars.block_512[16][2] ;
 wire \sha256cu.m_pad_pars.block_512[16][3] ;
 wire \sha256cu.m_pad_pars.block_512[16][4] ;
 wire \sha256cu.m_pad_pars.block_512[16][5] ;
 wire \sha256cu.m_pad_pars.block_512[16][6] ;
 wire \sha256cu.m_pad_pars.block_512[16][7] ;
 wire \sha256cu.m_pad_pars.block_512[17][0] ;
 wire \sha256cu.m_pad_pars.block_512[17][1] ;
 wire \sha256cu.m_pad_pars.block_512[17][2] ;
 wire \sha256cu.m_pad_pars.block_512[17][3] ;
 wire \sha256cu.m_pad_pars.block_512[17][4] ;
 wire \sha256cu.m_pad_pars.block_512[17][5] ;
 wire \sha256cu.m_pad_pars.block_512[17][6] ;
 wire \sha256cu.m_pad_pars.block_512[17][7] ;
 wire \sha256cu.m_pad_pars.block_512[18][0] ;
 wire \sha256cu.m_pad_pars.block_512[18][1] ;
 wire \sha256cu.m_pad_pars.block_512[18][2] ;
 wire \sha256cu.m_pad_pars.block_512[18][3] ;
 wire \sha256cu.m_pad_pars.block_512[18][4] ;
 wire \sha256cu.m_pad_pars.block_512[18][5] ;
 wire \sha256cu.m_pad_pars.block_512[18][6] ;
 wire \sha256cu.m_pad_pars.block_512[18][7] ;
 wire \sha256cu.m_pad_pars.block_512[19][0] ;
 wire \sha256cu.m_pad_pars.block_512[19][1] ;
 wire \sha256cu.m_pad_pars.block_512[19][2] ;
 wire \sha256cu.m_pad_pars.block_512[19][3] ;
 wire \sha256cu.m_pad_pars.block_512[19][4] ;
 wire \sha256cu.m_pad_pars.block_512[19][5] ;
 wire \sha256cu.m_pad_pars.block_512[19][6] ;
 wire \sha256cu.m_pad_pars.block_512[19][7] ;
 wire \sha256cu.m_pad_pars.block_512[1][0] ;
 wire \sha256cu.m_pad_pars.block_512[1][1] ;
 wire \sha256cu.m_pad_pars.block_512[1][2] ;
 wire \sha256cu.m_pad_pars.block_512[1][3] ;
 wire \sha256cu.m_pad_pars.block_512[1][4] ;
 wire \sha256cu.m_pad_pars.block_512[1][5] ;
 wire \sha256cu.m_pad_pars.block_512[1][6] ;
 wire \sha256cu.m_pad_pars.block_512[1][7] ;
 wire \sha256cu.m_pad_pars.block_512[20][0] ;
 wire \sha256cu.m_pad_pars.block_512[20][1] ;
 wire \sha256cu.m_pad_pars.block_512[20][2] ;
 wire \sha256cu.m_pad_pars.block_512[20][3] ;
 wire \sha256cu.m_pad_pars.block_512[20][4] ;
 wire \sha256cu.m_pad_pars.block_512[20][5] ;
 wire \sha256cu.m_pad_pars.block_512[20][6] ;
 wire \sha256cu.m_pad_pars.block_512[20][7] ;
 wire \sha256cu.m_pad_pars.block_512[21][0] ;
 wire \sha256cu.m_pad_pars.block_512[21][1] ;
 wire \sha256cu.m_pad_pars.block_512[21][2] ;
 wire \sha256cu.m_pad_pars.block_512[21][3] ;
 wire \sha256cu.m_pad_pars.block_512[21][4] ;
 wire \sha256cu.m_pad_pars.block_512[21][5] ;
 wire \sha256cu.m_pad_pars.block_512[21][6] ;
 wire \sha256cu.m_pad_pars.block_512[21][7] ;
 wire \sha256cu.m_pad_pars.block_512[22][0] ;
 wire \sha256cu.m_pad_pars.block_512[22][1] ;
 wire \sha256cu.m_pad_pars.block_512[22][2] ;
 wire \sha256cu.m_pad_pars.block_512[22][3] ;
 wire \sha256cu.m_pad_pars.block_512[22][4] ;
 wire \sha256cu.m_pad_pars.block_512[22][5] ;
 wire \sha256cu.m_pad_pars.block_512[22][6] ;
 wire \sha256cu.m_pad_pars.block_512[22][7] ;
 wire \sha256cu.m_pad_pars.block_512[23][0] ;
 wire \sha256cu.m_pad_pars.block_512[23][1] ;
 wire \sha256cu.m_pad_pars.block_512[23][2] ;
 wire \sha256cu.m_pad_pars.block_512[23][3] ;
 wire \sha256cu.m_pad_pars.block_512[23][4] ;
 wire \sha256cu.m_pad_pars.block_512[23][5] ;
 wire \sha256cu.m_pad_pars.block_512[23][6] ;
 wire \sha256cu.m_pad_pars.block_512[23][7] ;
 wire \sha256cu.m_pad_pars.block_512[24][0] ;
 wire \sha256cu.m_pad_pars.block_512[24][1] ;
 wire \sha256cu.m_pad_pars.block_512[24][2] ;
 wire \sha256cu.m_pad_pars.block_512[24][3] ;
 wire \sha256cu.m_pad_pars.block_512[24][4] ;
 wire \sha256cu.m_pad_pars.block_512[24][5] ;
 wire \sha256cu.m_pad_pars.block_512[24][6] ;
 wire \sha256cu.m_pad_pars.block_512[24][7] ;
 wire \sha256cu.m_pad_pars.block_512[25][0] ;
 wire \sha256cu.m_pad_pars.block_512[25][1] ;
 wire \sha256cu.m_pad_pars.block_512[25][2] ;
 wire \sha256cu.m_pad_pars.block_512[25][3] ;
 wire \sha256cu.m_pad_pars.block_512[25][4] ;
 wire \sha256cu.m_pad_pars.block_512[25][5] ;
 wire \sha256cu.m_pad_pars.block_512[25][6] ;
 wire \sha256cu.m_pad_pars.block_512[25][7] ;
 wire \sha256cu.m_pad_pars.block_512[26][0] ;
 wire \sha256cu.m_pad_pars.block_512[26][1] ;
 wire \sha256cu.m_pad_pars.block_512[26][2] ;
 wire \sha256cu.m_pad_pars.block_512[26][3] ;
 wire \sha256cu.m_pad_pars.block_512[26][4] ;
 wire \sha256cu.m_pad_pars.block_512[26][5] ;
 wire \sha256cu.m_pad_pars.block_512[26][6] ;
 wire \sha256cu.m_pad_pars.block_512[26][7] ;
 wire \sha256cu.m_pad_pars.block_512[27][0] ;
 wire \sha256cu.m_pad_pars.block_512[27][1] ;
 wire \sha256cu.m_pad_pars.block_512[27][2] ;
 wire \sha256cu.m_pad_pars.block_512[27][3] ;
 wire \sha256cu.m_pad_pars.block_512[27][4] ;
 wire \sha256cu.m_pad_pars.block_512[27][5] ;
 wire \sha256cu.m_pad_pars.block_512[27][6] ;
 wire \sha256cu.m_pad_pars.block_512[27][7] ;
 wire \sha256cu.m_pad_pars.block_512[28][0] ;
 wire \sha256cu.m_pad_pars.block_512[28][1] ;
 wire \sha256cu.m_pad_pars.block_512[28][2] ;
 wire \sha256cu.m_pad_pars.block_512[28][3] ;
 wire \sha256cu.m_pad_pars.block_512[28][4] ;
 wire \sha256cu.m_pad_pars.block_512[28][5] ;
 wire \sha256cu.m_pad_pars.block_512[28][6] ;
 wire \sha256cu.m_pad_pars.block_512[28][7] ;
 wire \sha256cu.m_pad_pars.block_512[29][0] ;
 wire \sha256cu.m_pad_pars.block_512[29][1] ;
 wire \sha256cu.m_pad_pars.block_512[29][2] ;
 wire \sha256cu.m_pad_pars.block_512[29][3] ;
 wire \sha256cu.m_pad_pars.block_512[29][4] ;
 wire \sha256cu.m_pad_pars.block_512[29][5] ;
 wire \sha256cu.m_pad_pars.block_512[29][6] ;
 wire \sha256cu.m_pad_pars.block_512[29][7] ;
 wire \sha256cu.m_pad_pars.block_512[2][0] ;
 wire \sha256cu.m_pad_pars.block_512[2][1] ;
 wire \sha256cu.m_pad_pars.block_512[2][2] ;
 wire \sha256cu.m_pad_pars.block_512[2][3] ;
 wire \sha256cu.m_pad_pars.block_512[2][4] ;
 wire \sha256cu.m_pad_pars.block_512[2][5] ;
 wire \sha256cu.m_pad_pars.block_512[2][6] ;
 wire \sha256cu.m_pad_pars.block_512[2][7] ;
 wire \sha256cu.m_pad_pars.block_512[30][0] ;
 wire \sha256cu.m_pad_pars.block_512[30][1] ;
 wire \sha256cu.m_pad_pars.block_512[30][2] ;
 wire \sha256cu.m_pad_pars.block_512[30][3] ;
 wire \sha256cu.m_pad_pars.block_512[30][4] ;
 wire \sha256cu.m_pad_pars.block_512[30][5] ;
 wire \sha256cu.m_pad_pars.block_512[30][6] ;
 wire \sha256cu.m_pad_pars.block_512[30][7] ;
 wire \sha256cu.m_pad_pars.block_512[31][0] ;
 wire \sha256cu.m_pad_pars.block_512[31][1] ;
 wire \sha256cu.m_pad_pars.block_512[31][2] ;
 wire \sha256cu.m_pad_pars.block_512[31][3] ;
 wire \sha256cu.m_pad_pars.block_512[31][4] ;
 wire \sha256cu.m_pad_pars.block_512[31][5] ;
 wire \sha256cu.m_pad_pars.block_512[31][6] ;
 wire \sha256cu.m_pad_pars.block_512[31][7] ;
 wire \sha256cu.m_pad_pars.block_512[32][0] ;
 wire \sha256cu.m_pad_pars.block_512[32][1] ;
 wire \sha256cu.m_pad_pars.block_512[32][2] ;
 wire \sha256cu.m_pad_pars.block_512[32][3] ;
 wire \sha256cu.m_pad_pars.block_512[32][4] ;
 wire \sha256cu.m_pad_pars.block_512[32][5] ;
 wire \sha256cu.m_pad_pars.block_512[32][6] ;
 wire \sha256cu.m_pad_pars.block_512[32][7] ;
 wire \sha256cu.m_pad_pars.block_512[33][0] ;
 wire \sha256cu.m_pad_pars.block_512[33][1] ;
 wire \sha256cu.m_pad_pars.block_512[33][2] ;
 wire \sha256cu.m_pad_pars.block_512[33][3] ;
 wire \sha256cu.m_pad_pars.block_512[33][4] ;
 wire \sha256cu.m_pad_pars.block_512[33][5] ;
 wire \sha256cu.m_pad_pars.block_512[33][6] ;
 wire \sha256cu.m_pad_pars.block_512[33][7] ;
 wire \sha256cu.m_pad_pars.block_512[34][0] ;
 wire \sha256cu.m_pad_pars.block_512[34][1] ;
 wire \sha256cu.m_pad_pars.block_512[34][2] ;
 wire \sha256cu.m_pad_pars.block_512[34][3] ;
 wire \sha256cu.m_pad_pars.block_512[34][4] ;
 wire \sha256cu.m_pad_pars.block_512[34][5] ;
 wire \sha256cu.m_pad_pars.block_512[34][6] ;
 wire \sha256cu.m_pad_pars.block_512[34][7] ;
 wire \sha256cu.m_pad_pars.block_512[35][0] ;
 wire \sha256cu.m_pad_pars.block_512[35][1] ;
 wire \sha256cu.m_pad_pars.block_512[35][2] ;
 wire \sha256cu.m_pad_pars.block_512[35][3] ;
 wire \sha256cu.m_pad_pars.block_512[35][4] ;
 wire \sha256cu.m_pad_pars.block_512[35][5] ;
 wire \sha256cu.m_pad_pars.block_512[35][6] ;
 wire \sha256cu.m_pad_pars.block_512[35][7] ;
 wire \sha256cu.m_pad_pars.block_512[36][0] ;
 wire \sha256cu.m_pad_pars.block_512[36][1] ;
 wire \sha256cu.m_pad_pars.block_512[36][2] ;
 wire \sha256cu.m_pad_pars.block_512[36][3] ;
 wire \sha256cu.m_pad_pars.block_512[36][4] ;
 wire \sha256cu.m_pad_pars.block_512[36][5] ;
 wire \sha256cu.m_pad_pars.block_512[36][6] ;
 wire \sha256cu.m_pad_pars.block_512[36][7] ;
 wire \sha256cu.m_pad_pars.block_512[37][0] ;
 wire \sha256cu.m_pad_pars.block_512[37][1] ;
 wire \sha256cu.m_pad_pars.block_512[37][2] ;
 wire \sha256cu.m_pad_pars.block_512[37][3] ;
 wire \sha256cu.m_pad_pars.block_512[37][4] ;
 wire \sha256cu.m_pad_pars.block_512[37][5] ;
 wire \sha256cu.m_pad_pars.block_512[37][6] ;
 wire \sha256cu.m_pad_pars.block_512[37][7] ;
 wire \sha256cu.m_pad_pars.block_512[38][0] ;
 wire \sha256cu.m_pad_pars.block_512[38][1] ;
 wire \sha256cu.m_pad_pars.block_512[38][2] ;
 wire \sha256cu.m_pad_pars.block_512[38][3] ;
 wire \sha256cu.m_pad_pars.block_512[38][4] ;
 wire \sha256cu.m_pad_pars.block_512[38][5] ;
 wire \sha256cu.m_pad_pars.block_512[38][6] ;
 wire \sha256cu.m_pad_pars.block_512[38][7] ;
 wire \sha256cu.m_pad_pars.block_512[39][0] ;
 wire \sha256cu.m_pad_pars.block_512[39][1] ;
 wire \sha256cu.m_pad_pars.block_512[39][2] ;
 wire \sha256cu.m_pad_pars.block_512[39][3] ;
 wire \sha256cu.m_pad_pars.block_512[39][4] ;
 wire \sha256cu.m_pad_pars.block_512[39][5] ;
 wire \sha256cu.m_pad_pars.block_512[39][6] ;
 wire \sha256cu.m_pad_pars.block_512[39][7] ;
 wire \sha256cu.m_pad_pars.block_512[3][0] ;
 wire \sha256cu.m_pad_pars.block_512[3][1] ;
 wire \sha256cu.m_pad_pars.block_512[3][2] ;
 wire \sha256cu.m_pad_pars.block_512[3][3] ;
 wire \sha256cu.m_pad_pars.block_512[3][4] ;
 wire \sha256cu.m_pad_pars.block_512[3][5] ;
 wire \sha256cu.m_pad_pars.block_512[3][6] ;
 wire \sha256cu.m_pad_pars.block_512[3][7] ;
 wire \sha256cu.m_pad_pars.block_512[40][0] ;
 wire \sha256cu.m_pad_pars.block_512[40][1] ;
 wire \sha256cu.m_pad_pars.block_512[40][2] ;
 wire \sha256cu.m_pad_pars.block_512[40][3] ;
 wire \sha256cu.m_pad_pars.block_512[40][4] ;
 wire \sha256cu.m_pad_pars.block_512[40][5] ;
 wire \sha256cu.m_pad_pars.block_512[40][6] ;
 wire \sha256cu.m_pad_pars.block_512[40][7] ;
 wire \sha256cu.m_pad_pars.block_512[41][0] ;
 wire \sha256cu.m_pad_pars.block_512[41][1] ;
 wire \sha256cu.m_pad_pars.block_512[41][2] ;
 wire \sha256cu.m_pad_pars.block_512[41][3] ;
 wire \sha256cu.m_pad_pars.block_512[41][4] ;
 wire \sha256cu.m_pad_pars.block_512[41][5] ;
 wire \sha256cu.m_pad_pars.block_512[41][6] ;
 wire \sha256cu.m_pad_pars.block_512[41][7] ;
 wire \sha256cu.m_pad_pars.block_512[42][0] ;
 wire \sha256cu.m_pad_pars.block_512[42][1] ;
 wire \sha256cu.m_pad_pars.block_512[42][2] ;
 wire \sha256cu.m_pad_pars.block_512[42][3] ;
 wire \sha256cu.m_pad_pars.block_512[42][4] ;
 wire \sha256cu.m_pad_pars.block_512[42][5] ;
 wire \sha256cu.m_pad_pars.block_512[42][6] ;
 wire \sha256cu.m_pad_pars.block_512[42][7] ;
 wire \sha256cu.m_pad_pars.block_512[43][0] ;
 wire \sha256cu.m_pad_pars.block_512[43][1] ;
 wire \sha256cu.m_pad_pars.block_512[43][2] ;
 wire \sha256cu.m_pad_pars.block_512[43][3] ;
 wire \sha256cu.m_pad_pars.block_512[43][4] ;
 wire \sha256cu.m_pad_pars.block_512[43][5] ;
 wire \sha256cu.m_pad_pars.block_512[43][6] ;
 wire \sha256cu.m_pad_pars.block_512[43][7] ;
 wire \sha256cu.m_pad_pars.block_512[44][0] ;
 wire \sha256cu.m_pad_pars.block_512[44][1] ;
 wire \sha256cu.m_pad_pars.block_512[44][2] ;
 wire \sha256cu.m_pad_pars.block_512[44][3] ;
 wire \sha256cu.m_pad_pars.block_512[44][4] ;
 wire \sha256cu.m_pad_pars.block_512[44][5] ;
 wire \sha256cu.m_pad_pars.block_512[44][6] ;
 wire \sha256cu.m_pad_pars.block_512[44][7] ;
 wire \sha256cu.m_pad_pars.block_512[45][0] ;
 wire \sha256cu.m_pad_pars.block_512[45][1] ;
 wire \sha256cu.m_pad_pars.block_512[45][2] ;
 wire \sha256cu.m_pad_pars.block_512[45][3] ;
 wire \sha256cu.m_pad_pars.block_512[45][4] ;
 wire \sha256cu.m_pad_pars.block_512[45][5] ;
 wire \sha256cu.m_pad_pars.block_512[45][6] ;
 wire \sha256cu.m_pad_pars.block_512[45][7] ;
 wire \sha256cu.m_pad_pars.block_512[46][0] ;
 wire \sha256cu.m_pad_pars.block_512[46][1] ;
 wire \sha256cu.m_pad_pars.block_512[46][2] ;
 wire \sha256cu.m_pad_pars.block_512[46][3] ;
 wire \sha256cu.m_pad_pars.block_512[46][4] ;
 wire \sha256cu.m_pad_pars.block_512[46][5] ;
 wire \sha256cu.m_pad_pars.block_512[46][6] ;
 wire \sha256cu.m_pad_pars.block_512[46][7] ;
 wire \sha256cu.m_pad_pars.block_512[47][0] ;
 wire \sha256cu.m_pad_pars.block_512[47][1] ;
 wire \sha256cu.m_pad_pars.block_512[47][2] ;
 wire \sha256cu.m_pad_pars.block_512[47][3] ;
 wire \sha256cu.m_pad_pars.block_512[47][4] ;
 wire \sha256cu.m_pad_pars.block_512[47][5] ;
 wire \sha256cu.m_pad_pars.block_512[47][6] ;
 wire \sha256cu.m_pad_pars.block_512[47][7] ;
 wire \sha256cu.m_pad_pars.block_512[48][0] ;
 wire \sha256cu.m_pad_pars.block_512[48][1] ;
 wire \sha256cu.m_pad_pars.block_512[48][2] ;
 wire \sha256cu.m_pad_pars.block_512[48][3] ;
 wire \sha256cu.m_pad_pars.block_512[48][4] ;
 wire \sha256cu.m_pad_pars.block_512[48][5] ;
 wire \sha256cu.m_pad_pars.block_512[48][6] ;
 wire \sha256cu.m_pad_pars.block_512[48][7] ;
 wire \sha256cu.m_pad_pars.block_512[49][0] ;
 wire \sha256cu.m_pad_pars.block_512[49][1] ;
 wire \sha256cu.m_pad_pars.block_512[49][2] ;
 wire \sha256cu.m_pad_pars.block_512[49][3] ;
 wire \sha256cu.m_pad_pars.block_512[49][4] ;
 wire \sha256cu.m_pad_pars.block_512[49][5] ;
 wire \sha256cu.m_pad_pars.block_512[49][6] ;
 wire \sha256cu.m_pad_pars.block_512[49][7] ;
 wire \sha256cu.m_pad_pars.block_512[4][0] ;
 wire \sha256cu.m_pad_pars.block_512[4][1] ;
 wire \sha256cu.m_pad_pars.block_512[4][2] ;
 wire \sha256cu.m_pad_pars.block_512[4][3] ;
 wire \sha256cu.m_pad_pars.block_512[4][4] ;
 wire \sha256cu.m_pad_pars.block_512[4][5] ;
 wire \sha256cu.m_pad_pars.block_512[4][6] ;
 wire \sha256cu.m_pad_pars.block_512[4][7] ;
 wire \sha256cu.m_pad_pars.block_512[50][0] ;
 wire \sha256cu.m_pad_pars.block_512[50][1] ;
 wire \sha256cu.m_pad_pars.block_512[50][2] ;
 wire \sha256cu.m_pad_pars.block_512[50][3] ;
 wire \sha256cu.m_pad_pars.block_512[50][4] ;
 wire \sha256cu.m_pad_pars.block_512[50][5] ;
 wire \sha256cu.m_pad_pars.block_512[50][6] ;
 wire \sha256cu.m_pad_pars.block_512[50][7] ;
 wire \sha256cu.m_pad_pars.block_512[51][0] ;
 wire \sha256cu.m_pad_pars.block_512[51][1] ;
 wire \sha256cu.m_pad_pars.block_512[51][2] ;
 wire \sha256cu.m_pad_pars.block_512[51][3] ;
 wire \sha256cu.m_pad_pars.block_512[51][4] ;
 wire \sha256cu.m_pad_pars.block_512[51][5] ;
 wire \sha256cu.m_pad_pars.block_512[51][6] ;
 wire \sha256cu.m_pad_pars.block_512[51][7] ;
 wire \sha256cu.m_pad_pars.block_512[52][0] ;
 wire \sha256cu.m_pad_pars.block_512[52][1] ;
 wire \sha256cu.m_pad_pars.block_512[52][2] ;
 wire \sha256cu.m_pad_pars.block_512[52][3] ;
 wire \sha256cu.m_pad_pars.block_512[52][4] ;
 wire \sha256cu.m_pad_pars.block_512[52][5] ;
 wire \sha256cu.m_pad_pars.block_512[52][6] ;
 wire \sha256cu.m_pad_pars.block_512[52][7] ;
 wire \sha256cu.m_pad_pars.block_512[53][0] ;
 wire \sha256cu.m_pad_pars.block_512[53][1] ;
 wire \sha256cu.m_pad_pars.block_512[53][2] ;
 wire \sha256cu.m_pad_pars.block_512[53][3] ;
 wire \sha256cu.m_pad_pars.block_512[53][4] ;
 wire \sha256cu.m_pad_pars.block_512[53][5] ;
 wire \sha256cu.m_pad_pars.block_512[53][6] ;
 wire \sha256cu.m_pad_pars.block_512[53][7] ;
 wire \sha256cu.m_pad_pars.block_512[54][0] ;
 wire \sha256cu.m_pad_pars.block_512[54][1] ;
 wire \sha256cu.m_pad_pars.block_512[54][2] ;
 wire \sha256cu.m_pad_pars.block_512[54][3] ;
 wire \sha256cu.m_pad_pars.block_512[54][4] ;
 wire \sha256cu.m_pad_pars.block_512[54][5] ;
 wire \sha256cu.m_pad_pars.block_512[54][6] ;
 wire \sha256cu.m_pad_pars.block_512[54][7] ;
 wire \sha256cu.m_pad_pars.block_512[55][0] ;
 wire \sha256cu.m_pad_pars.block_512[55][1] ;
 wire \sha256cu.m_pad_pars.block_512[55][2] ;
 wire \sha256cu.m_pad_pars.block_512[55][3] ;
 wire \sha256cu.m_pad_pars.block_512[55][4] ;
 wire \sha256cu.m_pad_pars.block_512[55][5] ;
 wire \sha256cu.m_pad_pars.block_512[55][6] ;
 wire \sha256cu.m_pad_pars.block_512[55][7] ;
 wire \sha256cu.m_pad_pars.block_512[56][0] ;
 wire \sha256cu.m_pad_pars.block_512[56][1] ;
 wire \sha256cu.m_pad_pars.block_512[56][2] ;
 wire \sha256cu.m_pad_pars.block_512[56][3] ;
 wire \sha256cu.m_pad_pars.block_512[56][4] ;
 wire \sha256cu.m_pad_pars.block_512[56][5] ;
 wire \sha256cu.m_pad_pars.block_512[56][6] ;
 wire \sha256cu.m_pad_pars.block_512[56][7] ;
 wire \sha256cu.m_pad_pars.block_512[57][0] ;
 wire \sha256cu.m_pad_pars.block_512[57][1] ;
 wire \sha256cu.m_pad_pars.block_512[57][2] ;
 wire \sha256cu.m_pad_pars.block_512[57][3] ;
 wire \sha256cu.m_pad_pars.block_512[57][4] ;
 wire \sha256cu.m_pad_pars.block_512[57][5] ;
 wire \sha256cu.m_pad_pars.block_512[57][6] ;
 wire \sha256cu.m_pad_pars.block_512[57][7] ;
 wire \sha256cu.m_pad_pars.block_512[58][0] ;
 wire \sha256cu.m_pad_pars.block_512[58][1] ;
 wire \sha256cu.m_pad_pars.block_512[58][2] ;
 wire \sha256cu.m_pad_pars.block_512[58][3] ;
 wire \sha256cu.m_pad_pars.block_512[58][4] ;
 wire \sha256cu.m_pad_pars.block_512[58][5] ;
 wire \sha256cu.m_pad_pars.block_512[58][6] ;
 wire \sha256cu.m_pad_pars.block_512[58][7] ;
 wire \sha256cu.m_pad_pars.block_512[59][0] ;
 wire \sha256cu.m_pad_pars.block_512[59][1] ;
 wire \sha256cu.m_pad_pars.block_512[59][2] ;
 wire \sha256cu.m_pad_pars.block_512[59][3] ;
 wire \sha256cu.m_pad_pars.block_512[59][4] ;
 wire \sha256cu.m_pad_pars.block_512[59][5] ;
 wire \sha256cu.m_pad_pars.block_512[59][6] ;
 wire \sha256cu.m_pad_pars.block_512[59][7] ;
 wire \sha256cu.m_pad_pars.block_512[5][0] ;
 wire \sha256cu.m_pad_pars.block_512[5][1] ;
 wire \sha256cu.m_pad_pars.block_512[5][2] ;
 wire \sha256cu.m_pad_pars.block_512[5][3] ;
 wire \sha256cu.m_pad_pars.block_512[5][4] ;
 wire \sha256cu.m_pad_pars.block_512[5][5] ;
 wire \sha256cu.m_pad_pars.block_512[5][6] ;
 wire \sha256cu.m_pad_pars.block_512[5][7] ;
 wire \sha256cu.m_pad_pars.block_512[60][0] ;
 wire \sha256cu.m_pad_pars.block_512[60][1] ;
 wire \sha256cu.m_pad_pars.block_512[60][2] ;
 wire \sha256cu.m_pad_pars.block_512[60][3] ;
 wire \sha256cu.m_pad_pars.block_512[60][4] ;
 wire \sha256cu.m_pad_pars.block_512[60][5] ;
 wire \sha256cu.m_pad_pars.block_512[60][6] ;
 wire \sha256cu.m_pad_pars.block_512[60][7] ;
 wire \sha256cu.m_pad_pars.block_512[61][0] ;
 wire \sha256cu.m_pad_pars.block_512[61][1] ;
 wire \sha256cu.m_pad_pars.block_512[61][2] ;
 wire \sha256cu.m_pad_pars.block_512[61][3] ;
 wire \sha256cu.m_pad_pars.block_512[61][4] ;
 wire \sha256cu.m_pad_pars.block_512[61][5] ;
 wire \sha256cu.m_pad_pars.block_512[61][6] ;
 wire \sha256cu.m_pad_pars.block_512[61][7] ;
 wire \sha256cu.m_pad_pars.block_512[62][0] ;
 wire \sha256cu.m_pad_pars.block_512[62][1] ;
 wire \sha256cu.m_pad_pars.block_512[62][2] ;
 wire \sha256cu.m_pad_pars.block_512[62][3] ;
 wire \sha256cu.m_pad_pars.block_512[62][4] ;
 wire \sha256cu.m_pad_pars.block_512[62][5] ;
 wire \sha256cu.m_pad_pars.block_512[62][6] ;
 wire \sha256cu.m_pad_pars.block_512[62][7] ;
 wire \sha256cu.m_pad_pars.block_512[63][0] ;
 wire \sha256cu.m_pad_pars.block_512[63][1] ;
 wire \sha256cu.m_pad_pars.block_512[63][2] ;
 wire \sha256cu.m_pad_pars.block_512[63][3] ;
 wire \sha256cu.m_pad_pars.block_512[63][4] ;
 wire \sha256cu.m_pad_pars.block_512[63][5] ;
 wire \sha256cu.m_pad_pars.block_512[63][6] ;
 wire \sha256cu.m_pad_pars.block_512[63][7] ;
 wire \sha256cu.m_pad_pars.block_512[6][0] ;
 wire \sha256cu.m_pad_pars.block_512[6][1] ;
 wire \sha256cu.m_pad_pars.block_512[6][2] ;
 wire \sha256cu.m_pad_pars.block_512[6][3] ;
 wire \sha256cu.m_pad_pars.block_512[6][4] ;
 wire \sha256cu.m_pad_pars.block_512[6][5] ;
 wire \sha256cu.m_pad_pars.block_512[6][6] ;
 wire \sha256cu.m_pad_pars.block_512[6][7] ;
 wire \sha256cu.m_pad_pars.block_512[7][0] ;
 wire \sha256cu.m_pad_pars.block_512[7][1] ;
 wire \sha256cu.m_pad_pars.block_512[7][2] ;
 wire \sha256cu.m_pad_pars.block_512[7][3] ;
 wire \sha256cu.m_pad_pars.block_512[7][4] ;
 wire \sha256cu.m_pad_pars.block_512[7][5] ;
 wire \sha256cu.m_pad_pars.block_512[7][6] ;
 wire \sha256cu.m_pad_pars.block_512[7][7] ;
 wire \sha256cu.m_pad_pars.block_512[8][0] ;
 wire \sha256cu.m_pad_pars.block_512[8][1] ;
 wire \sha256cu.m_pad_pars.block_512[8][2] ;
 wire \sha256cu.m_pad_pars.block_512[8][3] ;
 wire \sha256cu.m_pad_pars.block_512[8][4] ;
 wire \sha256cu.m_pad_pars.block_512[8][5] ;
 wire \sha256cu.m_pad_pars.block_512[8][6] ;
 wire \sha256cu.m_pad_pars.block_512[8][7] ;
 wire \sha256cu.m_pad_pars.block_512[9][0] ;
 wire \sha256cu.m_pad_pars.block_512[9][1] ;
 wire \sha256cu.m_pad_pars.block_512[9][2] ;
 wire \sha256cu.m_pad_pars.block_512[9][3] ;
 wire \sha256cu.m_pad_pars.block_512[9][4] ;
 wire \sha256cu.m_pad_pars.block_512[9][5] ;
 wire \sha256cu.m_pad_pars.block_512[9][6] ;
 wire \sha256cu.m_pad_pars.block_512[9][7] ;
 wire \sha256cu.m_pad_pars.m_size[3] ;
 wire \sha256cu.m_pad_pars.m_size[4] ;
 wire \sha256cu.m_pad_pars.m_size[5] ;
 wire \sha256cu.m_pad_pars.m_size[6] ;
 wire \sha256cu.m_pad_pars.m_size[7] ;
 wire \sha256cu.m_pad_pars.m_size[8] ;
 wire \sha256cu.m_pad_pars.m_size[9] ;
 wire \sha256cu.m_pad_pars.temp_chk ;
 wire \sha256cu.msg_scheduler.counter_iteration[0] ;
 wire \sha256cu.msg_scheduler.counter_iteration[1] ;
 wire \sha256cu.msg_scheduler.counter_iteration[2] ;
 wire \sha256cu.msg_scheduler.counter_iteration[3] ;
 wire \sha256cu.msg_scheduler.counter_iteration[4] ;
 wire \sha256cu.msg_scheduler.counter_iteration[5] ;
 wire \sha256cu.msg_scheduler.counter_iteration[6] ;
 wire \sha256cu.msg_scheduler.mreg_0[0] ;
 wire \sha256cu.msg_scheduler.mreg_0[10] ;
 wire \sha256cu.msg_scheduler.mreg_0[11] ;
 wire \sha256cu.msg_scheduler.mreg_0[12] ;
 wire \sha256cu.msg_scheduler.mreg_0[13] ;
 wire \sha256cu.msg_scheduler.mreg_0[14] ;
 wire \sha256cu.msg_scheduler.mreg_0[15] ;
 wire \sha256cu.msg_scheduler.mreg_0[16] ;
 wire \sha256cu.msg_scheduler.mreg_0[17] ;
 wire \sha256cu.msg_scheduler.mreg_0[18] ;
 wire \sha256cu.msg_scheduler.mreg_0[19] ;
 wire \sha256cu.msg_scheduler.mreg_0[1] ;
 wire \sha256cu.msg_scheduler.mreg_0[20] ;
 wire \sha256cu.msg_scheduler.mreg_0[21] ;
 wire \sha256cu.msg_scheduler.mreg_0[22] ;
 wire \sha256cu.msg_scheduler.mreg_0[23] ;
 wire \sha256cu.msg_scheduler.mreg_0[24] ;
 wire \sha256cu.msg_scheduler.mreg_0[25] ;
 wire \sha256cu.msg_scheduler.mreg_0[26] ;
 wire \sha256cu.msg_scheduler.mreg_0[27] ;
 wire \sha256cu.msg_scheduler.mreg_0[28] ;
 wire \sha256cu.msg_scheduler.mreg_0[29] ;
 wire \sha256cu.msg_scheduler.mreg_0[2] ;
 wire \sha256cu.msg_scheduler.mreg_0[30] ;
 wire \sha256cu.msg_scheduler.mreg_0[31] ;
 wire \sha256cu.msg_scheduler.mreg_0[3] ;
 wire \sha256cu.msg_scheduler.mreg_0[4] ;
 wire \sha256cu.msg_scheduler.mreg_0[5] ;
 wire \sha256cu.msg_scheduler.mreg_0[6] ;
 wire \sha256cu.msg_scheduler.mreg_0[7] ;
 wire \sha256cu.msg_scheduler.mreg_0[8] ;
 wire \sha256cu.msg_scheduler.mreg_0[9] ;
 wire \sha256cu.msg_scheduler.mreg_10[0] ;
 wire \sha256cu.msg_scheduler.mreg_10[10] ;
 wire \sha256cu.msg_scheduler.mreg_10[11] ;
 wire \sha256cu.msg_scheduler.mreg_10[12] ;
 wire \sha256cu.msg_scheduler.mreg_10[13] ;
 wire \sha256cu.msg_scheduler.mreg_10[14] ;
 wire \sha256cu.msg_scheduler.mreg_10[15] ;
 wire \sha256cu.msg_scheduler.mreg_10[16] ;
 wire \sha256cu.msg_scheduler.mreg_10[17] ;
 wire \sha256cu.msg_scheduler.mreg_10[18] ;
 wire \sha256cu.msg_scheduler.mreg_10[19] ;
 wire \sha256cu.msg_scheduler.mreg_10[1] ;
 wire \sha256cu.msg_scheduler.mreg_10[20] ;
 wire \sha256cu.msg_scheduler.mreg_10[21] ;
 wire \sha256cu.msg_scheduler.mreg_10[22] ;
 wire \sha256cu.msg_scheduler.mreg_10[23] ;
 wire \sha256cu.msg_scheduler.mreg_10[24] ;
 wire \sha256cu.msg_scheduler.mreg_10[25] ;
 wire \sha256cu.msg_scheduler.mreg_10[26] ;
 wire \sha256cu.msg_scheduler.mreg_10[27] ;
 wire \sha256cu.msg_scheduler.mreg_10[28] ;
 wire \sha256cu.msg_scheduler.mreg_10[29] ;
 wire \sha256cu.msg_scheduler.mreg_10[2] ;
 wire \sha256cu.msg_scheduler.mreg_10[30] ;
 wire \sha256cu.msg_scheduler.mreg_10[31] ;
 wire \sha256cu.msg_scheduler.mreg_10[3] ;
 wire \sha256cu.msg_scheduler.mreg_10[4] ;
 wire \sha256cu.msg_scheduler.mreg_10[5] ;
 wire \sha256cu.msg_scheduler.mreg_10[6] ;
 wire \sha256cu.msg_scheduler.mreg_10[7] ;
 wire \sha256cu.msg_scheduler.mreg_10[8] ;
 wire \sha256cu.msg_scheduler.mreg_10[9] ;
 wire \sha256cu.msg_scheduler.mreg_11[0] ;
 wire \sha256cu.msg_scheduler.mreg_11[10] ;
 wire \sha256cu.msg_scheduler.mreg_11[11] ;
 wire \sha256cu.msg_scheduler.mreg_11[12] ;
 wire \sha256cu.msg_scheduler.mreg_11[13] ;
 wire \sha256cu.msg_scheduler.mreg_11[14] ;
 wire \sha256cu.msg_scheduler.mreg_11[15] ;
 wire \sha256cu.msg_scheduler.mreg_11[16] ;
 wire \sha256cu.msg_scheduler.mreg_11[17] ;
 wire \sha256cu.msg_scheduler.mreg_11[18] ;
 wire \sha256cu.msg_scheduler.mreg_11[19] ;
 wire \sha256cu.msg_scheduler.mreg_11[1] ;
 wire \sha256cu.msg_scheduler.mreg_11[20] ;
 wire \sha256cu.msg_scheduler.mreg_11[21] ;
 wire \sha256cu.msg_scheduler.mreg_11[22] ;
 wire \sha256cu.msg_scheduler.mreg_11[23] ;
 wire \sha256cu.msg_scheduler.mreg_11[24] ;
 wire \sha256cu.msg_scheduler.mreg_11[25] ;
 wire \sha256cu.msg_scheduler.mreg_11[26] ;
 wire \sha256cu.msg_scheduler.mreg_11[27] ;
 wire \sha256cu.msg_scheduler.mreg_11[28] ;
 wire \sha256cu.msg_scheduler.mreg_11[29] ;
 wire \sha256cu.msg_scheduler.mreg_11[2] ;
 wire \sha256cu.msg_scheduler.mreg_11[30] ;
 wire \sha256cu.msg_scheduler.mreg_11[31] ;
 wire \sha256cu.msg_scheduler.mreg_11[3] ;
 wire \sha256cu.msg_scheduler.mreg_11[4] ;
 wire \sha256cu.msg_scheduler.mreg_11[5] ;
 wire \sha256cu.msg_scheduler.mreg_11[6] ;
 wire \sha256cu.msg_scheduler.mreg_11[7] ;
 wire \sha256cu.msg_scheduler.mreg_11[8] ;
 wire \sha256cu.msg_scheduler.mreg_11[9] ;
 wire \sha256cu.msg_scheduler.mreg_12[0] ;
 wire \sha256cu.msg_scheduler.mreg_12[10] ;
 wire \sha256cu.msg_scheduler.mreg_12[11] ;
 wire \sha256cu.msg_scheduler.mreg_12[12] ;
 wire \sha256cu.msg_scheduler.mreg_12[13] ;
 wire \sha256cu.msg_scheduler.mreg_12[14] ;
 wire \sha256cu.msg_scheduler.mreg_12[15] ;
 wire \sha256cu.msg_scheduler.mreg_12[16] ;
 wire \sha256cu.msg_scheduler.mreg_12[17] ;
 wire \sha256cu.msg_scheduler.mreg_12[18] ;
 wire \sha256cu.msg_scheduler.mreg_12[19] ;
 wire \sha256cu.msg_scheduler.mreg_12[1] ;
 wire \sha256cu.msg_scheduler.mreg_12[20] ;
 wire \sha256cu.msg_scheduler.mreg_12[21] ;
 wire \sha256cu.msg_scheduler.mreg_12[22] ;
 wire \sha256cu.msg_scheduler.mreg_12[23] ;
 wire \sha256cu.msg_scheduler.mreg_12[24] ;
 wire \sha256cu.msg_scheduler.mreg_12[25] ;
 wire \sha256cu.msg_scheduler.mreg_12[26] ;
 wire \sha256cu.msg_scheduler.mreg_12[27] ;
 wire \sha256cu.msg_scheduler.mreg_12[28] ;
 wire \sha256cu.msg_scheduler.mreg_12[29] ;
 wire \sha256cu.msg_scheduler.mreg_12[2] ;
 wire \sha256cu.msg_scheduler.mreg_12[30] ;
 wire \sha256cu.msg_scheduler.mreg_12[31] ;
 wire \sha256cu.msg_scheduler.mreg_12[3] ;
 wire \sha256cu.msg_scheduler.mreg_12[4] ;
 wire \sha256cu.msg_scheduler.mreg_12[5] ;
 wire \sha256cu.msg_scheduler.mreg_12[6] ;
 wire \sha256cu.msg_scheduler.mreg_12[7] ;
 wire \sha256cu.msg_scheduler.mreg_12[8] ;
 wire \sha256cu.msg_scheduler.mreg_12[9] ;
 wire \sha256cu.msg_scheduler.mreg_13[0] ;
 wire \sha256cu.msg_scheduler.mreg_13[10] ;
 wire \sha256cu.msg_scheduler.mreg_13[11] ;
 wire \sha256cu.msg_scheduler.mreg_13[12] ;
 wire \sha256cu.msg_scheduler.mreg_13[13] ;
 wire \sha256cu.msg_scheduler.mreg_13[14] ;
 wire \sha256cu.msg_scheduler.mreg_13[15] ;
 wire \sha256cu.msg_scheduler.mreg_13[16] ;
 wire \sha256cu.msg_scheduler.mreg_13[17] ;
 wire \sha256cu.msg_scheduler.mreg_13[18] ;
 wire \sha256cu.msg_scheduler.mreg_13[19] ;
 wire \sha256cu.msg_scheduler.mreg_13[1] ;
 wire \sha256cu.msg_scheduler.mreg_13[20] ;
 wire \sha256cu.msg_scheduler.mreg_13[21] ;
 wire \sha256cu.msg_scheduler.mreg_13[22] ;
 wire \sha256cu.msg_scheduler.mreg_13[23] ;
 wire \sha256cu.msg_scheduler.mreg_13[24] ;
 wire \sha256cu.msg_scheduler.mreg_13[25] ;
 wire \sha256cu.msg_scheduler.mreg_13[26] ;
 wire \sha256cu.msg_scheduler.mreg_13[27] ;
 wire \sha256cu.msg_scheduler.mreg_13[28] ;
 wire \sha256cu.msg_scheduler.mreg_13[29] ;
 wire \sha256cu.msg_scheduler.mreg_13[2] ;
 wire \sha256cu.msg_scheduler.mreg_13[30] ;
 wire \sha256cu.msg_scheduler.mreg_13[31] ;
 wire \sha256cu.msg_scheduler.mreg_13[3] ;
 wire \sha256cu.msg_scheduler.mreg_13[4] ;
 wire \sha256cu.msg_scheduler.mreg_13[5] ;
 wire \sha256cu.msg_scheduler.mreg_13[6] ;
 wire \sha256cu.msg_scheduler.mreg_13[7] ;
 wire \sha256cu.msg_scheduler.mreg_13[8] ;
 wire \sha256cu.msg_scheduler.mreg_13[9] ;
 wire \sha256cu.msg_scheduler.mreg_14[0] ;
 wire \sha256cu.msg_scheduler.mreg_14[10] ;
 wire \sha256cu.msg_scheduler.mreg_14[11] ;
 wire \sha256cu.msg_scheduler.mreg_14[12] ;
 wire \sha256cu.msg_scheduler.mreg_14[13] ;
 wire \sha256cu.msg_scheduler.mreg_14[14] ;
 wire \sha256cu.msg_scheduler.mreg_14[15] ;
 wire \sha256cu.msg_scheduler.mreg_14[16] ;
 wire \sha256cu.msg_scheduler.mreg_14[17] ;
 wire \sha256cu.msg_scheduler.mreg_14[18] ;
 wire \sha256cu.msg_scheduler.mreg_14[19] ;
 wire \sha256cu.msg_scheduler.mreg_14[1] ;
 wire \sha256cu.msg_scheduler.mreg_14[20] ;
 wire \sha256cu.msg_scheduler.mreg_14[21] ;
 wire \sha256cu.msg_scheduler.mreg_14[22] ;
 wire \sha256cu.msg_scheduler.mreg_14[23] ;
 wire \sha256cu.msg_scheduler.mreg_14[24] ;
 wire \sha256cu.msg_scheduler.mreg_14[25] ;
 wire \sha256cu.msg_scheduler.mreg_14[26] ;
 wire \sha256cu.msg_scheduler.mreg_14[27] ;
 wire \sha256cu.msg_scheduler.mreg_14[28] ;
 wire \sha256cu.msg_scheduler.mreg_14[29] ;
 wire \sha256cu.msg_scheduler.mreg_14[2] ;
 wire \sha256cu.msg_scheduler.mreg_14[30] ;
 wire \sha256cu.msg_scheduler.mreg_14[31] ;
 wire \sha256cu.msg_scheduler.mreg_14[3] ;
 wire \sha256cu.msg_scheduler.mreg_14[4] ;
 wire \sha256cu.msg_scheduler.mreg_14[5] ;
 wire \sha256cu.msg_scheduler.mreg_14[6] ;
 wire \sha256cu.msg_scheduler.mreg_14[7] ;
 wire \sha256cu.msg_scheduler.mreg_14[8] ;
 wire \sha256cu.msg_scheduler.mreg_14[9] ;
 wire \sha256cu.msg_scheduler.mreg_1[0] ;
 wire \sha256cu.msg_scheduler.mreg_1[10] ;
 wire \sha256cu.msg_scheduler.mreg_1[11] ;
 wire \sha256cu.msg_scheduler.mreg_1[12] ;
 wire \sha256cu.msg_scheduler.mreg_1[13] ;
 wire \sha256cu.msg_scheduler.mreg_1[14] ;
 wire \sha256cu.msg_scheduler.mreg_1[15] ;
 wire \sha256cu.msg_scheduler.mreg_1[16] ;
 wire \sha256cu.msg_scheduler.mreg_1[17] ;
 wire \sha256cu.msg_scheduler.mreg_1[18] ;
 wire \sha256cu.msg_scheduler.mreg_1[19] ;
 wire \sha256cu.msg_scheduler.mreg_1[1] ;
 wire \sha256cu.msg_scheduler.mreg_1[20] ;
 wire \sha256cu.msg_scheduler.mreg_1[21] ;
 wire \sha256cu.msg_scheduler.mreg_1[22] ;
 wire \sha256cu.msg_scheduler.mreg_1[23] ;
 wire \sha256cu.msg_scheduler.mreg_1[24] ;
 wire \sha256cu.msg_scheduler.mreg_1[25] ;
 wire \sha256cu.msg_scheduler.mreg_1[26] ;
 wire \sha256cu.msg_scheduler.mreg_1[27] ;
 wire \sha256cu.msg_scheduler.mreg_1[28] ;
 wire \sha256cu.msg_scheduler.mreg_1[29] ;
 wire \sha256cu.msg_scheduler.mreg_1[2] ;
 wire \sha256cu.msg_scheduler.mreg_1[30] ;
 wire \sha256cu.msg_scheduler.mreg_1[31] ;
 wire \sha256cu.msg_scheduler.mreg_1[3] ;
 wire \sha256cu.msg_scheduler.mreg_1[4] ;
 wire \sha256cu.msg_scheduler.mreg_1[5] ;
 wire \sha256cu.msg_scheduler.mreg_1[6] ;
 wire \sha256cu.msg_scheduler.mreg_1[7] ;
 wire \sha256cu.msg_scheduler.mreg_1[8] ;
 wire \sha256cu.msg_scheduler.mreg_1[9] ;
 wire \sha256cu.msg_scheduler.mreg_2[0] ;
 wire \sha256cu.msg_scheduler.mreg_2[10] ;
 wire \sha256cu.msg_scheduler.mreg_2[11] ;
 wire \sha256cu.msg_scheduler.mreg_2[12] ;
 wire \sha256cu.msg_scheduler.mreg_2[13] ;
 wire \sha256cu.msg_scheduler.mreg_2[14] ;
 wire \sha256cu.msg_scheduler.mreg_2[15] ;
 wire \sha256cu.msg_scheduler.mreg_2[16] ;
 wire \sha256cu.msg_scheduler.mreg_2[17] ;
 wire \sha256cu.msg_scheduler.mreg_2[18] ;
 wire \sha256cu.msg_scheduler.mreg_2[19] ;
 wire \sha256cu.msg_scheduler.mreg_2[1] ;
 wire \sha256cu.msg_scheduler.mreg_2[20] ;
 wire \sha256cu.msg_scheduler.mreg_2[21] ;
 wire \sha256cu.msg_scheduler.mreg_2[22] ;
 wire \sha256cu.msg_scheduler.mreg_2[23] ;
 wire \sha256cu.msg_scheduler.mreg_2[24] ;
 wire \sha256cu.msg_scheduler.mreg_2[25] ;
 wire \sha256cu.msg_scheduler.mreg_2[26] ;
 wire \sha256cu.msg_scheduler.mreg_2[27] ;
 wire \sha256cu.msg_scheduler.mreg_2[28] ;
 wire \sha256cu.msg_scheduler.mreg_2[29] ;
 wire \sha256cu.msg_scheduler.mreg_2[2] ;
 wire \sha256cu.msg_scheduler.mreg_2[30] ;
 wire \sha256cu.msg_scheduler.mreg_2[31] ;
 wire \sha256cu.msg_scheduler.mreg_2[3] ;
 wire \sha256cu.msg_scheduler.mreg_2[4] ;
 wire \sha256cu.msg_scheduler.mreg_2[5] ;
 wire \sha256cu.msg_scheduler.mreg_2[6] ;
 wire \sha256cu.msg_scheduler.mreg_2[7] ;
 wire \sha256cu.msg_scheduler.mreg_2[8] ;
 wire \sha256cu.msg_scheduler.mreg_2[9] ;
 wire \sha256cu.msg_scheduler.mreg_3[0] ;
 wire \sha256cu.msg_scheduler.mreg_3[10] ;
 wire \sha256cu.msg_scheduler.mreg_3[11] ;
 wire \sha256cu.msg_scheduler.mreg_3[12] ;
 wire \sha256cu.msg_scheduler.mreg_3[13] ;
 wire \sha256cu.msg_scheduler.mreg_3[14] ;
 wire \sha256cu.msg_scheduler.mreg_3[15] ;
 wire \sha256cu.msg_scheduler.mreg_3[16] ;
 wire \sha256cu.msg_scheduler.mreg_3[17] ;
 wire \sha256cu.msg_scheduler.mreg_3[18] ;
 wire \sha256cu.msg_scheduler.mreg_3[19] ;
 wire \sha256cu.msg_scheduler.mreg_3[1] ;
 wire \sha256cu.msg_scheduler.mreg_3[20] ;
 wire \sha256cu.msg_scheduler.mreg_3[21] ;
 wire \sha256cu.msg_scheduler.mreg_3[22] ;
 wire \sha256cu.msg_scheduler.mreg_3[23] ;
 wire \sha256cu.msg_scheduler.mreg_3[24] ;
 wire \sha256cu.msg_scheduler.mreg_3[25] ;
 wire \sha256cu.msg_scheduler.mreg_3[26] ;
 wire \sha256cu.msg_scheduler.mreg_3[27] ;
 wire \sha256cu.msg_scheduler.mreg_3[28] ;
 wire \sha256cu.msg_scheduler.mreg_3[29] ;
 wire \sha256cu.msg_scheduler.mreg_3[2] ;
 wire \sha256cu.msg_scheduler.mreg_3[30] ;
 wire \sha256cu.msg_scheduler.mreg_3[31] ;
 wire \sha256cu.msg_scheduler.mreg_3[3] ;
 wire \sha256cu.msg_scheduler.mreg_3[4] ;
 wire \sha256cu.msg_scheduler.mreg_3[5] ;
 wire \sha256cu.msg_scheduler.mreg_3[6] ;
 wire \sha256cu.msg_scheduler.mreg_3[7] ;
 wire \sha256cu.msg_scheduler.mreg_3[8] ;
 wire \sha256cu.msg_scheduler.mreg_3[9] ;
 wire \sha256cu.msg_scheduler.mreg_4[0] ;
 wire \sha256cu.msg_scheduler.mreg_4[10] ;
 wire \sha256cu.msg_scheduler.mreg_4[11] ;
 wire \sha256cu.msg_scheduler.mreg_4[12] ;
 wire \sha256cu.msg_scheduler.mreg_4[13] ;
 wire \sha256cu.msg_scheduler.mreg_4[14] ;
 wire \sha256cu.msg_scheduler.mreg_4[15] ;
 wire \sha256cu.msg_scheduler.mreg_4[16] ;
 wire \sha256cu.msg_scheduler.mreg_4[17] ;
 wire \sha256cu.msg_scheduler.mreg_4[18] ;
 wire \sha256cu.msg_scheduler.mreg_4[19] ;
 wire \sha256cu.msg_scheduler.mreg_4[1] ;
 wire \sha256cu.msg_scheduler.mreg_4[20] ;
 wire \sha256cu.msg_scheduler.mreg_4[21] ;
 wire \sha256cu.msg_scheduler.mreg_4[22] ;
 wire \sha256cu.msg_scheduler.mreg_4[23] ;
 wire \sha256cu.msg_scheduler.mreg_4[24] ;
 wire \sha256cu.msg_scheduler.mreg_4[25] ;
 wire \sha256cu.msg_scheduler.mreg_4[26] ;
 wire \sha256cu.msg_scheduler.mreg_4[27] ;
 wire \sha256cu.msg_scheduler.mreg_4[28] ;
 wire \sha256cu.msg_scheduler.mreg_4[29] ;
 wire \sha256cu.msg_scheduler.mreg_4[2] ;
 wire \sha256cu.msg_scheduler.mreg_4[30] ;
 wire \sha256cu.msg_scheduler.mreg_4[31] ;
 wire \sha256cu.msg_scheduler.mreg_4[3] ;
 wire \sha256cu.msg_scheduler.mreg_4[4] ;
 wire \sha256cu.msg_scheduler.mreg_4[5] ;
 wire \sha256cu.msg_scheduler.mreg_4[6] ;
 wire \sha256cu.msg_scheduler.mreg_4[7] ;
 wire \sha256cu.msg_scheduler.mreg_4[8] ;
 wire \sha256cu.msg_scheduler.mreg_4[9] ;
 wire \sha256cu.msg_scheduler.mreg_5[0] ;
 wire \sha256cu.msg_scheduler.mreg_5[10] ;
 wire \sha256cu.msg_scheduler.mreg_5[11] ;
 wire \sha256cu.msg_scheduler.mreg_5[12] ;
 wire \sha256cu.msg_scheduler.mreg_5[13] ;
 wire \sha256cu.msg_scheduler.mreg_5[14] ;
 wire \sha256cu.msg_scheduler.mreg_5[15] ;
 wire \sha256cu.msg_scheduler.mreg_5[16] ;
 wire \sha256cu.msg_scheduler.mreg_5[17] ;
 wire \sha256cu.msg_scheduler.mreg_5[18] ;
 wire \sha256cu.msg_scheduler.mreg_5[19] ;
 wire \sha256cu.msg_scheduler.mreg_5[1] ;
 wire \sha256cu.msg_scheduler.mreg_5[20] ;
 wire \sha256cu.msg_scheduler.mreg_5[21] ;
 wire \sha256cu.msg_scheduler.mreg_5[22] ;
 wire \sha256cu.msg_scheduler.mreg_5[23] ;
 wire \sha256cu.msg_scheduler.mreg_5[24] ;
 wire \sha256cu.msg_scheduler.mreg_5[25] ;
 wire \sha256cu.msg_scheduler.mreg_5[26] ;
 wire \sha256cu.msg_scheduler.mreg_5[27] ;
 wire \sha256cu.msg_scheduler.mreg_5[28] ;
 wire \sha256cu.msg_scheduler.mreg_5[29] ;
 wire \sha256cu.msg_scheduler.mreg_5[2] ;
 wire \sha256cu.msg_scheduler.mreg_5[30] ;
 wire \sha256cu.msg_scheduler.mreg_5[31] ;
 wire \sha256cu.msg_scheduler.mreg_5[3] ;
 wire \sha256cu.msg_scheduler.mreg_5[4] ;
 wire \sha256cu.msg_scheduler.mreg_5[5] ;
 wire \sha256cu.msg_scheduler.mreg_5[6] ;
 wire \sha256cu.msg_scheduler.mreg_5[7] ;
 wire \sha256cu.msg_scheduler.mreg_5[8] ;
 wire \sha256cu.msg_scheduler.mreg_5[9] ;
 wire \sha256cu.msg_scheduler.mreg_6[0] ;
 wire \sha256cu.msg_scheduler.mreg_6[10] ;
 wire \sha256cu.msg_scheduler.mreg_6[11] ;
 wire \sha256cu.msg_scheduler.mreg_6[12] ;
 wire \sha256cu.msg_scheduler.mreg_6[13] ;
 wire \sha256cu.msg_scheduler.mreg_6[14] ;
 wire \sha256cu.msg_scheduler.mreg_6[15] ;
 wire \sha256cu.msg_scheduler.mreg_6[16] ;
 wire \sha256cu.msg_scheduler.mreg_6[17] ;
 wire \sha256cu.msg_scheduler.mreg_6[18] ;
 wire \sha256cu.msg_scheduler.mreg_6[19] ;
 wire \sha256cu.msg_scheduler.mreg_6[1] ;
 wire \sha256cu.msg_scheduler.mreg_6[20] ;
 wire \sha256cu.msg_scheduler.mreg_6[21] ;
 wire \sha256cu.msg_scheduler.mreg_6[22] ;
 wire \sha256cu.msg_scheduler.mreg_6[23] ;
 wire \sha256cu.msg_scheduler.mreg_6[24] ;
 wire \sha256cu.msg_scheduler.mreg_6[25] ;
 wire \sha256cu.msg_scheduler.mreg_6[26] ;
 wire \sha256cu.msg_scheduler.mreg_6[27] ;
 wire \sha256cu.msg_scheduler.mreg_6[28] ;
 wire \sha256cu.msg_scheduler.mreg_6[29] ;
 wire \sha256cu.msg_scheduler.mreg_6[2] ;
 wire \sha256cu.msg_scheduler.mreg_6[30] ;
 wire \sha256cu.msg_scheduler.mreg_6[31] ;
 wire \sha256cu.msg_scheduler.mreg_6[3] ;
 wire \sha256cu.msg_scheduler.mreg_6[4] ;
 wire \sha256cu.msg_scheduler.mreg_6[5] ;
 wire \sha256cu.msg_scheduler.mreg_6[6] ;
 wire \sha256cu.msg_scheduler.mreg_6[7] ;
 wire \sha256cu.msg_scheduler.mreg_6[8] ;
 wire \sha256cu.msg_scheduler.mreg_6[9] ;
 wire \sha256cu.msg_scheduler.mreg_7[0] ;
 wire \sha256cu.msg_scheduler.mreg_7[10] ;
 wire \sha256cu.msg_scheduler.mreg_7[11] ;
 wire \sha256cu.msg_scheduler.mreg_7[12] ;
 wire \sha256cu.msg_scheduler.mreg_7[13] ;
 wire \sha256cu.msg_scheduler.mreg_7[14] ;
 wire \sha256cu.msg_scheduler.mreg_7[15] ;
 wire \sha256cu.msg_scheduler.mreg_7[16] ;
 wire \sha256cu.msg_scheduler.mreg_7[17] ;
 wire \sha256cu.msg_scheduler.mreg_7[18] ;
 wire \sha256cu.msg_scheduler.mreg_7[19] ;
 wire \sha256cu.msg_scheduler.mreg_7[1] ;
 wire \sha256cu.msg_scheduler.mreg_7[20] ;
 wire \sha256cu.msg_scheduler.mreg_7[21] ;
 wire \sha256cu.msg_scheduler.mreg_7[22] ;
 wire \sha256cu.msg_scheduler.mreg_7[23] ;
 wire \sha256cu.msg_scheduler.mreg_7[24] ;
 wire \sha256cu.msg_scheduler.mreg_7[25] ;
 wire \sha256cu.msg_scheduler.mreg_7[26] ;
 wire \sha256cu.msg_scheduler.mreg_7[27] ;
 wire \sha256cu.msg_scheduler.mreg_7[28] ;
 wire \sha256cu.msg_scheduler.mreg_7[29] ;
 wire \sha256cu.msg_scheduler.mreg_7[2] ;
 wire \sha256cu.msg_scheduler.mreg_7[30] ;
 wire \sha256cu.msg_scheduler.mreg_7[31] ;
 wire \sha256cu.msg_scheduler.mreg_7[3] ;
 wire \sha256cu.msg_scheduler.mreg_7[4] ;
 wire \sha256cu.msg_scheduler.mreg_7[5] ;
 wire \sha256cu.msg_scheduler.mreg_7[6] ;
 wire \sha256cu.msg_scheduler.mreg_7[7] ;
 wire \sha256cu.msg_scheduler.mreg_7[8] ;
 wire \sha256cu.msg_scheduler.mreg_7[9] ;
 wire \sha256cu.msg_scheduler.mreg_8[0] ;
 wire \sha256cu.msg_scheduler.mreg_8[10] ;
 wire \sha256cu.msg_scheduler.mreg_8[11] ;
 wire \sha256cu.msg_scheduler.mreg_8[12] ;
 wire \sha256cu.msg_scheduler.mreg_8[13] ;
 wire \sha256cu.msg_scheduler.mreg_8[14] ;
 wire \sha256cu.msg_scheduler.mreg_8[15] ;
 wire \sha256cu.msg_scheduler.mreg_8[16] ;
 wire \sha256cu.msg_scheduler.mreg_8[17] ;
 wire \sha256cu.msg_scheduler.mreg_8[18] ;
 wire \sha256cu.msg_scheduler.mreg_8[19] ;
 wire \sha256cu.msg_scheduler.mreg_8[1] ;
 wire \sha256cu.msg_scheduler.mreg_8[20] ;
 wire \sha256cu.msg_scheduler.mreg_8[21] ;
 wire \sha256cu.msg_scheduler.mreg_8[22] ;
 wire \sha256cu.msg_scheduler.mreg_8[23] ;
 wire \sha256cu.msg_scheduler.mreg_8[24] ;
 wire \sha256cu.msg_scheduler.mreg_8[25] ;
 wire \sha256cu.msg_scheduler.mreg_8[26] ;
 wire \sha256cu.msg_scheduler.mreg_8[27] ;
 wire \sha256cu.msg_scheduler.mreg_8[28] ;
 wire \sha256cu.msg_scheduler.mreg_8[29] ;
 wire \sha256cu.msg_scheduler.mreg_8[2] ;
 wire \sha256cu.msg_scheduler.mreg_8[30] ;
 wire \sha256cu.msg_scheduler.mreg_8[31] ;
 wire \sha256cu.msg_scheduler.mreg_8[3] ;
 wire \sha256cu.msg_scheduler.mreg_8[4] ;
 wire \sha256cu.msg_scheduler.mreg_8[5] ;
 wire \sha256cu.msg_scheduler.mreg_8[6] ;
 wire \sha256cu.msg_scheduler.mreg_8[7] ;
 wire \sha256cu.msg_scheduler.mreg_8[8] ;
 wire \sha256cu.msg_scheduler.mreg_8[9] ;
 wire \sha256cu.msg_scheduler.mreg_9[0] ;
 wire \sha256cu.msg_scheduler.mreg_9[10] ;
 wire \sha256cu.msg_scheduler.mreg_9[11] ;
 wire \sha256cu.msg_scheduler.mreg_9[12] ;
 wire \sha256cu.msg_scheduler.mreg_9[13] ;
 wire \sha256cu.msg_scheduler.mreg_9[14] ;
 wire \sha256cu.msg_scheduler.mreg_9[15] ;
 wire \sha256cu.msg_scheduler.mreg_9[16] ;
 wire \sha256cu.msg_scheduler.mreg_9[17] ;
 wire \sha256cu.msg_scheduler.mreg_9[18] ;
 wire \sha256cu.msg_scheduler.mreg_9[19] ;
 wire \sha256cu.msg_scheduler.mreg_9[1] ;
 wire \sha256cu.msg_scheduler.mreg_9[20] ;
 wire \sha256cu.msg_scheduler.mreg_9[21] ;
 wire \sha256cu.msg_scheduler.mreg_9[22] ;
 wire \sha256cu.msg_scheduler.mreg_9[23] ;
 wire \sha256cu.msg_scheduler.mreg_9[24] ;
 wire \sha256cu.msg_scheduler.mreg_9[25] ;
 wire \sha256cu.msg_scheduler.mreg_9[26] ;
 wire \sha256cu.msg_scheduler.mreg_9[27] ;
 wire \sha256cu.msg_scheduler.mreg_9[28] ;
 wire \sha256cu.msg_scheduler.mreg_9[29] ;
 wire \sha256cu.msg_scheduler.mreg_9[2] ;
 wire \sha256cu.msg_scheduler.mreg_9[30] ;
 wire \sha256cu.msg_scheduler.mreg_9[31] ;
 wire \sha256cu.msg_scheduler.mreg_9[3] ;
 wire \sha256cu.msg_scheduler.mreg_9[4] ;
 wire \sha256cu.msg_scheduler.mreg_9[5] ;
 wire \sha256cu.msg_scheduler.mreg_9[6] ;
 wire \sha256cu.msg_scheduler.mreg_9[7] ;
 wire \sha256cu.msg_scheduler.mreg_9[8] ;
 wire \sha256cu.msg_scheduler.mreg_9[9] ;
 wire \sha256cu.msg_scheduler.temp_case ;
 wire \sha256cu.temp_case ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__or2_1 _06775_ (.A(net257),
    .B(\state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01474_));
 sky130_fd_sc_hd__clkbuf_1 _06776_ (.A(_01474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00032_));
 sky130_fd_sc_hd__or4_2 _06777_ (.A(net201),
    .B(net234),
    .C(net223),
    .D(net256),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01475_));
 sky130_fd_sc_hd__or4_2 _06778_ (.A(net112),
    .B(net190),
    .C(net179),
    .D(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01476_));
 sky130_fd_sc_hd__or4_1 _06779_ (.A(net34),
    .B(net67),
    .C(net56),
    .D(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01477_));
 sky130_fd_sc_hd__or4_2 _06780_ (.A(net245),
    .B(net23),
    .C(net12),
    .D(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01478_));
 sky130_fd_sc_hd__or4_4 _06781_ (.A(net78),
    .B(net111),
    .C(net100),
    .D(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01479_));
 sky130_fd_sc_hd__or4_2 _06782_ (.A(net123),
    .B(net156),
    .C(net145),
    .D(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01480_));
 sky130_fd_sc_hd__or4_1 _06783_ (.A(_01477_),
    .B(_01478_),
    .C(_01479_),
    .D(_01480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01481_));
 sky130_fd_sc_hd__or4_1 _06784_ (.A(net195),
    .B(net198),
    .C(net197),
    .D(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01482_));
 sky130_fd_sc_hd__or4_4 _06785_ (.A(net191),
    .B(net194),
    .C(net193),
    .D(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01483_));
 sky130_fd_sc_hd__or4_2 _06786_ (.A(net199),
    .B(net203),
    .C(net202),
    .D(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01484_));
 sky130_fd_sc_hd__or4_2 _06787_ (.A(net204),
    .B(net207),
    .C(net206),
    .D(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01485_));
 sky130_fd_sc_hd__or4_1 _06788_ (.A(_01482_),
    .B(_01483_),
    .C(_01484_),
    .D(_01485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01486_));
 sky130_fd_sc_hd__or4_2 _06789_ (.A(net177),
    .B(net181),
    .C(net180),
    .D(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01487_));
 sky130_fd_sc_hd__or4_1 _06790_ (.A(net167),
    .B(net176),
    .C(net175),
    .D(net178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01488_));
 sky130_fd_sc_hd__or4_1 _06791_ (.A(net182),
    .B(net185),
    .C(net184),
    .D(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01489_));
 sky130_fd_sc_hd__or4_2 _06792_ (.A(net186),
    .B(net189),
    .C(net188),
    .D(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01490_));
 sky130_fd_sc_hd__or4_2 _06793_ (.A(_01487_),
    .B(_01488_),
    .C(_01489_),
    .D(_01490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01491_));
 sky130_fd_sc_hd__or4_2 _06794_ (.A(net213),
    .B(net216),
    .C(net215),
    .D(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01492_));
 sky130_fd_sc_hd__or4_2 _06795_ (.A(net208),
    .B(net211),
    .C(net210),
    .D(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01493_));
 sky130_fd_sc_hd__or4_2 _06796_ (.A(net217),
    .B(net220),
    .C(net219),
    .D(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01494_));
 sky130_fd_sc_hd__or4_2 _06797_ (.A(net221),
    .B(net225),
    .C(net224),
    .D(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01495_));
 sky130_fd_sc_hd__or4_1 _06798_ (.A(_01492_),
    .B(_01493_),
    .C(_01494_),
    .D(_01495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01496_));
 sky130_fd_sc_hd__or4_2 _06799_ (.A(net230),
    .B(net233),
    .C(net232),
    .D(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01497_));
 sky130_fd_sc_hd__or4_2 _06800_ (.A(net226),
    .B(net229),
    .C(net228),
    .D(net231),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01498_));
 sky130_fd_sc_hd__or4_1 _06801_ (.A(net235),
    .B(net238),
    .C(net237),
    .D(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01499_));
 sky130_fd_sc_hd__or4_1 _06802_ (.A(net239),
    .B(net242),
    .C(net241),
    .D(net244),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01500_));
 sky130_fd_sc_hd__or4_1 _06803_ (.A(_01497_),
    .B(_01498_),
    .C(_01499_),
    .D(_01500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01501_));
 sky130_fd_sc_hd__or4_1 _06804_ (.A(_01486_),
    .B(_01491_),
    .C(_01496_),
    .D(_01501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01502_));
 sky130_fd_sc_hd__or4_1 _06805_ (.A(_01475_),
    .B(_01476_),
    .C(_01481_),
    .D(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01503_));
 sky130_fd_sc_hd__xor2_1 _06806_ (.A(Hash_Digest),
    .B(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01504_));
 sky130_fd_sc_hd__or4_1 _06807_ (.A(net165),
    .B(net169),
    .C(net168),
    .D(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01505_));
 sky130_fd_sc_hd__or4_2 _06808_ (.A(net170),
    .B(net173),
    .C(net172),
    .D(_01505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01506_));
 sky130_fd_sc_hd__or4_1 _06809_ (.A(net135),
    .B(net138),
    .C(net137),
    .D(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01507_));
 sky130_fd_sc_hd__or4_1 _06810_ (.A(net130),
    .B(net133),
    .C(net132),
    .D(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01508_));
 sky130_fd_sc_hd__or4_1 _06811_ (.A(net139),
    .B(net142),
    .C(net141),
    .D(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01509_));
 sky130_fd_sc_hd__or4_4 _06812_ (.A(net143),
    .B(net147),
    .C(net146),
    .D(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01510_));
 sky130_fd_sc_hd__or4_1 _06813_ (.A(_01507_),
    .B(_01508_),
    .C(_01509_),
    .D(_01510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01511_));
 sky130_fd_sc_hd__or4_4 _06814_ (.A(net152),
    .B(net155),
    .C(net154),
    .D(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01512_));
 sky130_fd_sc_hd__or4_2 _06815_ (.A(net148),
    .B(net151),
    .C(net150),
    .D(net153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01513_));
 sky130_fd_sc_hd__or4_2 _06816_ (.A(net157),
    .B(net160),
    .C(net159),
    .D(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01514_));
 sky130_fd_sc_hd__or4_1 _06817_ (.A(net161),
    .B(net164),
    .C(net163),
    .D(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01515_));
 sky130_fd_sc_hd__or4_1 _06818_ (.A(_01512_),
    .B(_01513_),
    .C(_01514_),
    .D(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01516_));
 sky130_fd_sc_hd__or4_1 _06819_ (.A(_01504_),
    .B(_01506_),
    .C(_01511_),
    .D(_01516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01517_));
 sky130_fd_sc_hd__or4_1 _06820_ (.A(net81),
    .B(net84),
    .C(net83),
    .D(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01518_));
 sky130_fd_sc_hd__or4_1 _06821_ (.A(net76),
    .B(net80),
    .C(net79),
    .D(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01519_));
 sky130_fd_sc_hd__or4_1 _06822_ (.A(net85),
    .B(net88),
    .C(net87),
    .D(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01520_));
 sky130_fd_sc_hd__or4_2 _06823_ (.A(net90),
    .B(net93),
    .C(net92),
    .D(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01521_));
 sky130_fd_sc_hd__or4_1 _06824_ (.A(_01518_),
    .B(_01519_),
    .C(_01520_),
    .D(_01521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01522_));
 sky130_fd_sc_hd__or4_4 _06825_ (.A(net63),
    .B(net66),
    .C(net65),
    .D(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01523_));
 sky130_fd_sc_hd__or4_2 _06826_ (.A(net59),
    .B(net62),
    .C(net61),
    .D(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01524_));
 sky130_fd_sc_hd__or4_1 _06827_ (.A(net68),
    .B(net71),
    .C(net70),
    .D(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01525_));
 sky130_fd_sc_hd__or4_2 _06828_ (.A(net72),
    .B(net75),
    .C(net74),
    .D(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01526_));
 sky130_fd_sc_hd__or4_1 _06829_ (.A(_01523_),
    .B(_01524_),
    .C(_01525_),
    .D(_01526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01527_));
 sky130_fd_sc_hd__or4_4 _06830_ (.A(net98),
    .B(net102),
    .C(net101),
    .D(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01528_));
 sky130_fd_sc_hd__or4_2 _06831_ (.A(net94),
    .B(net97),
    .C(net96),
    .D(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01529_));
 sky130_fd_sc_hd__or4_1 _06832_ (.A(net103),
    .B(net106),
    .C(net105),
    .D(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01530_));
 sky130_fd_sc_hd__or4_1 _06833_ (.A(net107),
    .B(net110),
    .C(net109),
    .D(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01531_));
 sky130_fd_sc_hd__or4_1 _06834_ (.A(_01528_),
    .B(_01529_),
    .C(_01530_),
    .D(_01531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01532_));
 sky130_fd_sc_hd__or4_1 _06835_ (.A(net117),
    .B(net120),
    .C(net119),
    .D(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01533_));
 sky130_fd_sc_hd__or4_1 _06836_ (.A(net113),
    .B(net116),
    .C(net115),
    .D(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01534_));
 sky130_fd_sc_hd__or4_1 _06837_ (.A(net121),
    .B(net125),
    .C(net124),
    .D(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01535_));
 sky130_fd_sc_hd__or4_1 _06838_ (.A(net126),
    .B(net129),
    .C(net128),
    .D(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01536_));
 sky130_fd_sc_hd__or4_2 _06839_ (.A(_01533_),
    .B(_01534_),
    .C(_01535_),
    .D(_01536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01537_));
 sky130_fd_sc_hd__or4_1 _06840_ (.A(_01522_),
    .B(_01527_),
    .C(_01532_),
    .D(_01537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01538_));
 sky130_fd_sc_hd__or4_1 _06841_ (.A(net10),
    .B(net14),
    .C(net13),
    .D(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01539_));
 sky130_fd_sc_hd__or4_1 _06842_ (.A(net6),
    .B(net9),
    .C(net8),
    .D(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01540_));
 sky130_fd_sc_hd__or4_2 _06843_ (.A(net15),
    .B(net18),
    .C(net17),
    .D(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01541_));
 sky130_fd_sc_hd__or4_1 _06844_ (.A(net19),
    .B(net22),
    .C(net21),
    .D(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01542_));
 sky130_fd_sc_hd__or4_1 _06845_ (.A(_01539_),
    .B(_01540_),
    .C(_01541_),
    .D(_01542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01543_));
 sky130_fd_sc_hd__or4_1 _06846_ (.A(net248),
    .B(net251),
    .C(net250),
    .D(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01544_));
 sky130_fd_sc_hd__or4_2 _06847_ (.A(net243),
    .B(net247),
    .C(net246),
    .D(net249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01545_));
 sky130_fd_sc_hd__or4_1 _06848_ (.A(net252),
    .B(net255),
    .C(net254),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01546_));
 sky130_fd_sc_hd__or4_2 _06849_ (.A(net2),
    .B(net5),
    .C(net4),
    .D(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01547_));
 sky130_fd_sc_hd__or4_1 _06850_ (.A(_01544_),
    .B(_01545_),
    .C(_01546_),
    .D(_01547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01548_));
 sky130_fd_sc_hd__or4_2 _06851_ (.A(net28),
    .B(net31),
    .C(net30),
    .D(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01549_));
 sky130_fd_sc_hd__or4_4 _06852_ (.A(net24),
    .B(net27),
    .C(net26),
    .D(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01550_));
 sky130_fd_sc_hd__or4_2 _06853_ (.A(net32),
    .B(net36),
    .C(net35),
    .D(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01551_));
 sky130_fd_sc_hd__or4_4 _06854_ (.A(net37),
    .B(net40),
    .C(net39),
    .D(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01552_));
 sky130_fd_sc_hd__or4_1 _06855_ (.A(_01549_),
    .B(_01550_),
    .C(_01551_),
    .D(_01552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01553_));
 sky130_fd_sc_hd__or4_4 _06856_ (.A(net46),
    .B(net49),
    .C(net48),
    .D(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01554_));
 sky130_fd_sc_hd__or4_2 _06857_ (.A(net41),
    .B(net44),
    .C(net43),
    .D(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01555_));
 sky130_fd_sc_hd__or4_1 _06858_ (.A(net50),
    .B(net53),
    .C(net52),
    .D(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01556_));
 sky130_fd_sc_hd__or4_1 _06859_ (.A(net54),
    .B(net58),
    .C(net57),
    .D(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01557_));
 sky130_fd_sc_hd__or4_2 _06860_ (.A(_01554_),
    .B(_01555_),
    .C(_01556_),
    .D(_01557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01558_));
 sky130_fd_sc_hd__or4_1 _06861_ (.A(_01543_),
    .B(_01548_),
    .C(_01553_),
    .D(_01558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01559_));
 sky130_fd_sc_hd__nor4_1 _06862_ (.A(_01503_),
    .B(_01517_),
    .C(_01538_),
    .D(_01559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01560_));
 sky130_fd_sc_hd__and2b_1 _06863_ (.A_N(_01560_),
    .B(\sha256cu.hashing_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01561_));
 sky130_fd_sc_hd__nor3b_1 _06864_ (.A(net257),
    .B(_01561_),
    .C_N(\state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00033_));
 sky130_fd_sc_hd__inv_2 _06865_ (.A(\state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01562_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(\state[1] ),
    .B(_01561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01563_));
 sky130_fd_sc_hd__a21oi_1 _06867_ (.A1(_01562_),
    .A2(_01563_),
    .B1(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00034_));
 sky130_fd_sc_hd__o21ba_1 _06868_ (.A1(\state[3] ),
    .A2(\state[2] ),
    .B1_N(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00035_));
 sky130_fd_sc_hd__buf_8 _06869_ (.A(\sha256cu.iter_processing.rst ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01564_));
 sky130_fd_sc_hd__or4_2 _06870_ (.A(\sha256cu.msg_scheduler.counter_iteration[0] ),
    .B(\sha256cu.msg_scheduler.counter_iteration[3] ),
    .C(\sha256cu.msg_scheduler.counter_iteration[2] ),
    .D(\sha256cu.msg_scheduler.counter_iteration[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01565_));
 sky130_fd_sc_hd__nor3_4 _06871_ (.A(\sha256cu.msg_scheduler.counter_iteration[5] ),
    .B(\sha256cu.msg_scheduler.counter_iteration[4] ),
    .C(_01565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01566_));
 sky130_fd_sc_hd__and2_1 _06872_ (.A(\sha256cu.msg_scheduler.counter_iteration[6] ),
    .B(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01567_));
 sky130_fd_sc_hd__o21a_2 _06873_ (.A1(\sha256cu.msg_scheduler.temp_case ),
    .A2(_01567_),
    .B1(\sha256cu.iter_processing.padding_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _06874_ (.A0(\sha256cu.counter_iteration[5] ),
    .A1(\sha256cu.msg_scheduler.counter_iteration[5] ),
    .S(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01569_));
 sky130_fd_sc_hd__nand2_4 _06875_ (.A(_01564_),
    .B(_01569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01570_));
 sky130_fd_sc_hd__clkinv_2 _06876_ (.A(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01571_));
 sky130_fd_sc_hd__clkbuf_4 _06877_ (.A(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_2 _06878_ (.A0(\sha256cu.counter_iteration[2] ),
    .A1(\sha256cu.msg_scheduler.counter_iteration[2] ),
    .S(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01572_));
 sky130_fd_sc_hd__nand2_8 _06879_ (.A(\sha256cu.iter_processing.rst ),
    .B(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01573_));
 sky130_fd_sc_hd__o21ai_1 _06880_ (.A1(\sha256cu.msg_scheduler.temp_case ),
    .A2(_01567_),
    .B1(\sha256cu.iter_processing.padding_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01574_));
 sky130_fd_sc_hd__or2_1 _06881_ (.A(\sha256cu.counter_iteration[0] ),
    .B(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01575_));
 sky130_fd_sc_hd__o211a_1 _06882_ (.A1(\sha256cu.msg_scheduler.counter_iteration[0] ),
    .A2(_01574_),
    .B1(_01575_),
    .C1(\sha256cu.iter_processing.rst ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01576_));
 sky130_fd_sc_hd__buf_6 _06883_ (.A(_01576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01577_));
 sky130_fd_sc_hd__nand2_4 _06884_ (.A(_01573_),
    .B(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01578_));
 sky130_fd_sc_hd__mux2_2 _06885_ (.A0(\sha256cu.counter_iteration[1] ),
    .A1(\sha256cu.msg_scheduler.counter_iteration[1] ),
    .S(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01579_));
 sky130_fd_sc_hd__buf_4 _06886_ (.A(_01579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01580_));
 sky130_fd_sc_hd__nor2_1 _06887_ (.A(_01578_),
    .B(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01581_));
 sky130_fd_sc_hd__mux2_1 _06888_ (.A0(\sha256cu.counter_iteration[4] ),
    .A1(\sha256cu.msg_scheduler.counter_iteration[4] ),
    .S(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01582_));
 sky130_fd_sc_hd__nand2_4 _06889_ (.A(_01564_),
    .B(_01582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01583_));
 sky130_fd_sc_hd__clkbuf_4 _06890_ (.A(_01583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01584_));
 sky130_fd_sc_hd__clkbuf_4 _06891_ (.A(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01585_));
 sky130_fd_sc_hd__and2_1 _06892_ (.A(_01573_),
    .B(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _06893_ (.A0(\sha256cu.counter_iteration[3] ),
    .A1(\sha256cu.msg_scheduler.counter_iteration[3] ),
    .S(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01587_));
 sky130_fd_sc_hd__nand2_4 _06894_ (.A(_01564_),
    .B(_01587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01588_));
 sky130_fd_sc_hd__clkinv_2 _06895_ (.A(_01588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01589_));
 sky130_fd_sc_hd__buf_4 _06896_ (.A(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01590_));
 sky130_fd_sc_hd__nor2_2 _06897_ (.A(_01586_),
    .B(_01590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01591_));
 sky130_fd_sc_hd__clkinv_2 _06898_ (.A(_01573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_2 _06899_ (.A(_01592_),
    .B(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01593_));
 sky130_fd_sc_hd__clkbuf_4 _06900_ (.A(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00452_));
 sky130_fd_sc_hd__or2_2 _06901_ (.A(_01592_),
    .B(_00452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01594_));
 sky130_fd_sc_hd__and3_2 _06902_ (.A(_01593_),
    .B(_01590_),
    .C(_01594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01595_));
 sky130_fd_sc_hd__inv_2 _06903_ (.A(_01583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01596_));
 sky130_fd_sc_hd__nor2_1 _06904_ (.A(_01593_),
    .B(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01597_));
 sky130_fd_sc_hd__or2_2 _06905_ (.A(_01596_),
    .B(_01597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01598_));
 sky130_fd_sc_hd__o32a_1 _06906_ (.A1(_01581_),
    .A2(_01585_),
    .A3(_01591_),
    .B1(_01595_),
    .B2(_01598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01599_));
 sky130_fd_sc_hd__nand2_4 _06907_ (.A(\sha256cu.iter_processing.rst ),
    .B(_01579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01600_));
 sky130_fd_sc_hd__clkinv_2 _06908_ (.A(_01600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00453_));
 sky130_fd_sc_hd__nor2_2 _06909_ (.A(_01592_),
    .B(_00453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01601_));
 sky130_fd_sc_hd__clkbuf_4 _06910_ (.A(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01602_));
 sky130_fd_sc_hd__clkbuf_4 _06911_ (.A(_01602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01603_));
 sky130_fd_sc_hd__nor2_2 _06912_ (.A(_01601_),
    .B(_01603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01604_));
 sky130_fd_sc_hd__clkinv_2 _06913_ (.A(_01579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01605_));
 sky130_fd_sc_hd__nand2_4 _06914_ (.A(_01577_),
    .B(_01605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01606_));
 sky130_fd_sc_hd__buf_4 _06915_ (.A(_01573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01607_));
 sky130_fd_sc_hd__nor2_8 _06916_ (.A(_01577_),
    .B(_01600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_2 _06917_ (.A(_01607_),
    .B(_01608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_2 _06918_ (.A(_01606_),
    .B(_01609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01610_));
 sky130_fd_sc_hd__clkbuf_4 _06919_ (.A(_01592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00454_));
 sky130_fd_sc_hd__nor2_2 _06920_ (.A(_00454_),
    .B(_01600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01611_));
 sky130_fd_sc_hd__nand2_4 _06921_ (.A(_01592_),
    .B(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01612_));
 sky130_fd_sc_hd__nand2_1 _06922_ (.A(_01589_),
    .B(_01612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01613_));
 sky130_fd_sc_hd__or2_1 _06923_ (.A(_01586_),
    .B(_01613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01614_));
 sky130_fd_sc_hd__or2_2 _06924_ (.A(_01611_),
    .B(_01614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01615_));
 sky130_fd_sc_hd__inv_2 _06925_ (.A(_01615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01616_));
 sky130_fd_sc_hd__clkbuf_4 _06926_ (.A(_01583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01617_));
 sky130_fd_sc_hd__clkbuf_4 _06927_ (.A(_01617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01618_));
 sky130_fd_sc_hd__a211o_1 _06928_ (.A1(_01604_),
    .A2(_01610_),
    .B1(_01616_),
    .C1(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01619_));
 sky130_fd_sc_hd__clkbuf_4 _06929_ (.A(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01620_));
 sky130_fd_sc_hd__clkbuf_4 _06930_ (.A(_01620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01621_));
 sky130_fd_sc_hd__nor2_2 _06931_ (.A(_00454_),
    .B(_01608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _06932_ (.A(_01606_),
    .B(_01588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_1 _06933_ (.A(_01622_),
    .B(_01623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01624_));
 sky130_fd_sc_hd__or2_2 _06934_ (.A(_01573_),
    .B(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01625_));
 sky130_fd_sc_hd__nand2_2 _06935_ (.A(_01625_),
    .B(_01612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01626_));
 sky130_fd_sc_hd__or2_1 _06936_ (.A(_01588_),
    .B(_01626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01627_));
 sky130_fd_sc_hd__nor2_1 _06937_ (.A(_01581_),
    .B(_01627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01628_));
 sky130_fd_sc_hd__clkbuf_4 _06938_ (.A(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01629_));
 sky130_fd_sc_hd__o31a_1 _06939_ (.A1(_01621_),
    .A2(_01624_),
    .A3(_01628_),
    .B1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01630_));
 sky130_fd_sc_hd__a2bb2o_1 _06940_ (.A1_N(_00457_),
    .A2_N(_01599_),
    .B1(_01619_),
    .B2(_01630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00000_));
 sky130_fd_sc_hd__clkbuf_4 _06941_ (.A(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01631_));
 sky130_fd_sc_hd__nor2_4 _06942_ (.A(_01573_),
    .B(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01632_));
 sky130_fd_sc_hd__nor2_2 _06943_ (.A(_01573_),
    .B(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01633_));
 sky130_fd_sc_hd__nor2_4 _06944_ (.A(_01632_),
    .B(_01633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01634_));
 sky130_fd_sc_hd__nand2_1 _06945_ (.A(_01586_),
    .B(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01635_));
 sky130_fd_sc_hd__and3_1 _06946_ (.A(_01590_),
    .B(_01634_),
    .C(_01635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01636_));
 sky130_fd_sc_hd__or2_2 _06947_ (.A(_00452_),
    .B(_00453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01637_));
 sky130_fd_sc_hd__and3_1 _06948_ (.A(_01578_),
    .B(_01637_),
    .C(_01612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01638_));
 sky130_fd_sc_hd__buf_2 _06949_ (.A(_01588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01639_));
 sky130_fd_sc_hd__clkbuf_4 _06950_ (.A(_01639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01640_));
 sky130_fd_sc_hd__or2_1 _06951_ (.A(_01601_),
    .B(_01640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01641_));
 sky130_fd_sc_hd__nand2_2 _06952_ (.A(_01577_),
    .B(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01642_));
 sky130_fd_sc_hd__nand2_2 _06953_ (.A(_01573_),
    .B(_01642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01643_));
 sky130_fd_sc_hd__clkbuf_4 _06954_ (.A(_01620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01644_));
 sky130_fd_sc_hd__o221a_1 _06955_ (.A1(_01636_),
    .A2(_01638_),
    .B1(_01641_),
    .B2(_01643_),
    .C1(_01644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01645_));
 sky130_fd_sc_hd__clkbuf_4 _06956_ (.A(_01590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01646_));
 sky130_fd_sc_hd__clkbuf_4 _06957_ (.A(_01646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01647_));
 sky130_fd_sc_hd__nand2_4 _06958_ (.A(_01573_),
    .B(_01606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_2 _06959_ (.A(_01608_),
    .B(_01648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01649_));
 sky130_fd_sc_hd__buf_2 _06960_ (.A(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01650_));
 sky130_fd_sc_hd__o221a_1 _06961_ (.A1(_01578_),
    .A2(_01647_),
    .B1(_01613_),
    .B2(_01649_),
    .C1(_01650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01651_));
 sky130_fd_sc_hd__clkbuf_4 _06962_ (.A(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01652_));
 sky130_fd_sc_hd__clkbuf_4 _06963_ (.A(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00456_));
 sky130_fd_sc_hd__clkbuf_4 _06964_ (.A(_01639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01653_));
 sky130_fd_sc_hd__or2_1 _06965_ (.A(_01608_),
    .B(_01648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01654_));
 sky130_fd_sc_hd__and3_1 _06966_ (.A(_01654_),
    .B(_01590_),
    .C(_01634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01655_));
 sky130_fd_sc_hd__a31o_1 _06967_ (.A1(_01607_),
    .A2(_01642_),
    .A3(_01653_),
    .B1(_01655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01656_));
 sky130_fd_sc_hd__clkbuf_4 _06968_ (.A(_01586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01657_));
 sky130_fd_sc_hd__nor2_2 _06969_ (.A(_01607_),
    .B(_01605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01658_));
 sky130_fd_sc_hd__or2_2 _06970_ (.A(_01601_),
    .B(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01659_));
 sky130_fd_sc_hd__nor2_1 _06971_ (.A(_01586_),
    .B(_01588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_2 _06972_ (.A(_01660_),
    .B(_01634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01661_));
 sky130_fd_sc_hd__o311a_1 _06973_ (.A1(_01657_),
    .A2(_01658_),
    .A3(_01659_),
    .B1(_01661_),
    .C1(_01617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01662_));
 sky130_fd_sc_hd__clkbuf_4 _06974_ (.A(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01663_));
 sky130_fd_sc_hd__a211o_1 _06975_ (.A1(_00456_),
    .A2(_01656_),
    .B1(_01662_),
    .C1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01664_));
 sky130_fd_sc_hd__o31ai_1 _06976_ (.A1(_01631_),
    .A2(_01645_),
    .A3(_01651_),
    .B1(_01664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00011_));
 sky130_fd_sc_hd__or2_2 _06977_ (.A(_00452_),
    .B(_01600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01665_));
 sky130_fd_sc_hd__nand2_4 _06978_ (.A(_00454_),
    .B(_01665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01666_));
 sky130_fd_sc_hd__nor2_4 _06979_ (.A(_01577_),
    .B(_00453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01667_));
 sky130_fd_sc_hd__o21a_1 _06980_ (.A1(_01667_),
    .A2(_01634_),
    .B1(_01591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01668_));
 sky130_fd_sc_hd__a21oi_1 _06981_ (.A1(_01646_),
    .A2(_01666_),
    .B1(_01668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01669_));
 sky130_fd_sc_hd__nor2_1 _06982_ (.A(_01632_),
    .B(_01649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01670_));
 sky130_fd_sc_hd__xnor2_1 _06983_ (.A(_01670_),
    .B(_01661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01671_));
 sky130_fd_sc_hd__mux2_1 _06984_ (.A0(_01669_),
    .A1(_01671_),
    .S(_01620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01672_));
 sky130_fd_sc_hd__or2_2 _06985_ (.A(_01608_),
    .B(_01623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01673_));
 sky130_fd_sc_hd__and3_1 _06986_ (.A(_01578_),
    .B(_01606_),
    .C(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01674_));
 sky130_fd_sc_hd__nor2_1 _06987_ (.A(_01602_),
    .B(_01626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01675_));
 sky130_fd_sc_hd__o21a_1 _06988_ (.A1(_01674_),
    .A2(_01675_),
    .B1(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01676_));
 sky130_fd_sc_hd__a31o_1 _06989_ (.A1(_01617_),
    .A2(_01661_),
    .A3(_01673_),
    .B1(_01676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _06990_ (.A0(_01672_),
    .A1(_01677_),
    .S(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01678_));
 sky130_fd_sc_hd__clkbuf_1 _06991_ (.A(_01678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00022_));
 sky130_fd_sc_hd__clkbuf_4 _06992_ (.A(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01679_));
 sky130_fd_sc_hd__clkbuf_4 _06993_ (.A(_01603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00455_));
 sky130_fd_sc_hd__nand2_1 _06994_ (.A(_00454_),
    .B(_01637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01680_));
 sky130_fd_sc_hd__and2_1 _06995_ (.A(_01648_),
    .B(_01680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01681_));
 sky130_fd_sc_hd__nor2_4 _06996_ (.A(_01590_),
    .B(_01633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01682_));
 sky130_fd_sc_hd__a221o_1 _06997_ (.A1(_00455_),
    .A2(_01681_),
    .B1(_01682_),
    .B2(_00452_),
    .C1(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01683_));
 sky130_fd_sc_hd__nand2_1 _06998_ (.A(_00452_),
    .B(_01658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01684_));
 sky130_fd_sc_hd__and3_1 _06999_ (.A(_01607_),
    .B(_01600_),
    .C(_01602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01685_));
 sky130_fd_sc_hd__a211o_1 _07000_ (.A1(_01604_),
    .A2(_01684_),
    .B1(_01685_),
    .C1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01686_));
 sky130_fd_sc_hd__clkbuf_4 _07001_ (.A(_01640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01687_));
 sky130_fd_sc_hd__nor2_1 _07002_ (.A(_01654_),
    .B(_01687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01688_));
 sky130_fd_sc_hd__nor2_2 _07003_ (.A(_00453_),
    .B(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01689_));
 sky130_fd_sc_hd__buf_2 _07004_ (.A(_01606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01690_));
 sky130_fd_sc_hd__or3_1 _07005_ (.A(_01583_),
    .B(_01597_),
    .C(_01689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01691_));
 sky130_fd_sc_hd__a31o_1 _07006_ (.A1(_01690_),
    .A2(_01603_),
    .A3(_01612_),
    .B1(_01691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01692_));
 sky130_fd_sc_hd__o311a_1 _07007_ (.A1(_01644_),
    .A2(_01688_),
    .A3(_01689_),
    .B1(_01692_),
    .C1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01693_));
 sky130_fd_sc_hd__a31o_1 _07008_ (.A1(_01679_),
    .A2(_01683_),
    .A3(_01686_),
    .B1(_01693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00025_));
 sky130_fd_sc_hd__nor2_2 _07009_ (.A(_01607_),
    .B(_01667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _07010_ (.A(_01640_),
    .B(_01694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01695_));
 sky130_fd_sc_hd__nor2_2 _07011_ (.A(_01667_),
    .B(_01634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01696_));
 sky130_fd_sc_hd__or3_1 _07012_ (.A(_01657_),
    .B(_01639_),
    .C(_01696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01697_));
 sky130_fd_sc_hd__inv_2 _07013_ (.A(_01691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01698_));
 sky130_fd_sc_hd__a32o_1 _07014_ (.A1(_01617_),
    .A2(_01614_),
    .A3(_01695_),
    .B1(_01697_),
    .B2(_01698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01699_));
 sky130_fd_sc_hd__nor2_1 _07015_ (.A(_01646_),
    .B(_01680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01700_));
 sky130_fd_sc_hd__nand2_2 _07016_ (.A(_01625_),
    .B(_01643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01701_));
 sky130_fd_sc_hd__inv_2 _07017_ (.A(_01626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01702_));
 sky130_fd_sc_hd__nor2_4 _07018_ (.A(_01601_),
    .B(_01588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(_01702_),
    .B(_01703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01704_));
 sky130_fd_sc_hd__o21ai_4 _07020_ (.A1(_01701_),
    .A2(_01704_),
    .B1(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_4 _07021_ (.A(_01607_),
    .B(_01608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01706_));
 sky130_fd_sc_hd__a31o_1 _07022_ (.A1(_01690_),
    .A2(_01640_),
    .A3(_01706_),
    .B1(_01595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01707_));
 sky130_fd_sc_hd__o22a_1 _07023_ (.A1(_01700_),
    .A2(_01705_),
    .B1(_01707_),
    .B2(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _07024_ (.A0(_01699_),
    .A1(_01708_),
    .S(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01709_));
 sky130_fd_sc_hd__clkbuf_1 _07025_ (.A(_01709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00026_));
 sky130_fd_sc_hd__nand2_1 _07026_ (.A(_01593_),
    .B(_01654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01710_));
 sky130_fd_sc_hd__nor2_1 _07027_ (.A(_01710_),
    .B(_01687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01711_));
 sky130_fd_sc_hd__nor2_1 _07028_ (.A(_01655_),
    .B(_01689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01712_));
 sky130_fd_sc_hd__o32a_1 _07029_ (.A1(_01598_),
    .A2(_01689_),
    .A3(_01711_),
    .B1(_01712_),
    .B2(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01713_));
 sky130_fd_sc_hd__and3_1 _07030_ (.A(_01606_),
    .B(_01602_),
    .C(_01706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01714_));
 sky130_fd_sc_hd__and3_1 _07031_ (.A(_01643_),
    .B(_01639_),
    .C(_01680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01715_));
 sky130_fd_sc_hd__a21o_1 _07032_ (.A1(_01666_),
    .A2(_01714_),
    .B1(_01715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01716_));
 sky130_fd_sc_hd__a21oi_1 _07033_ (.A1(_01682_),
    .A2(_01706_),
    .B1(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01717_));
 sky130_fd_sc_hd__a221o_1 _07034_ (.A1(_00456_),
    .A2(_01716_),
    .B1(_01717_),
    .B2(_01661_),
    .C1(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01718_));
 sky130_fd_sc_hd__o21a_1 _07035_ (.A1(_01679_),
    .A2(_01713_),
    .B1(_01718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00027_));
 sky130_fd_sc_hd__nand2_2 _07036_ (.A(_01578_),
    .B(_01625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01719_));
 sky130_fd_sc_hd__a22o_1 _07037_ (.A1(_01640_),
    .A2(_01719_),
    .B1(_01703_),
    .B2(_01690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01720_));
 sky130_fd_sc_hd__nor2_2 _07038_ (.A(_01667_),
    .B(_01590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01721_));
 sky130_fd_sc_hd__inv_2 _07039_ (.A(_01721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _07040_ (.A(_01602_),
    .B(_01684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01723_));
 sky130_fd_sc_hd__a21oi_1 _07041_ (.A1(_01722_),
    .A2(_01723_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01724_));
 sky130_fd_sc_hd__a21o_1 _07042_ (.A1(_01617_),
    .A2(_01720_),
    .B1(_01724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01725_));
 sky130_fd_sc_hd__o21ai_2 _07043_ (.A1(_00452_),
    .A2(_01590_),
    .B1(_01583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01726_));
 sky130_fd_sc_hd__nand2_1 _07044_ (.A(_01580_),
    .B(_01590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01727_));
 sky130_fd_sc_hd__nor2_1 _07045_ (.A(_00454_),
    .B(_01727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01728_));
 sky130_fd_sc_hd__a31o_1 _07046_ (.A1(_01607_),
    .A2(_01606_),
    .A3(_01588_),
    .B1(_01583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01729_));
 sky130_fd_sc_hd__o32a_1 _07047_ (.A1(_01609_),
    .A2(_01726_),
    .A3(_01728_),
    .B1(_01655_),
    .B2(_01729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01730_));
 sky130_fd_sc_hd__inv_2 _07048_ (.A(_01730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01731_));
 sky130_fd_sc_hd__mux2_1 _07049_ (.A0(_01725_),
    .A1(_01731_),
    .S(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01732_));
 sky130_fd_sc_hd__clkbuf_1 _07050_ (.A(_01732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _07051_ (.A(_01607_),
    .B(_01606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01733_));
 sky130_fd_sc_hd__o21ai_1 _07052_ (.A1(_01667_),
    .A2(_01614_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01734_));
 sky130_fd_sc_hd__a31o_1 _07053_ (.A1(_01648_),
    .A2(_01687_),
    .A3(_01733_),
    .B1(_01734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01735_));
 sky130_fd_sc_hd__o21ai_1 _07054_ (.A1(_01636_),
    .A2(_01689_),
    .B1(_00456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01736_));
 sky130_fd_sc_hd__o31a_1 _07055_ (.A1(_01657_),
    .A2(_01653_),
    .A3(_01611_),
    .B1(_01642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01737_));
 sky130_fd_sc_hd__nor2_1 _07056_ (.A(_01642_),
    .B(_01639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _07057_ (.A(_01690_),
    .B(_01666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01739_));
 sky130_fd_sc_hd__or3b_1 _07058_ (.A(_01726_),
    .B(_01739_),
    .C_N(_01706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01740_));
 sky130_fd_sc_hd__o311a_1 _07059_ (.A1(_01585_),
    .A2(_01737_),
    .A3(_01738_),
    .B1(_01740_),
    .C1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01741_));
 sky130_fd_sc_hd__a31o_1 _07060_ (.A1(_00457_),
    .A2(_01735_),
    .A3(_01736_),
    .B1(_01741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00029_));
 sky130_fd_sc_hd__a211o_1 _07061_ (.A1(_00455_),
    .A2(_01670_),
    .B1(_01675_),
    .C1(_00456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01742_));
 sky130_fd_sc_hd__or2_1 _07062_ (.A(_01667_),
    .B(_01643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01743_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(_01743_),
    .B(_01646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _07064_ (.A(_01626_),
    .B(_01744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01745_));
 sky130_fd_sc_hd__a311o_1 _07065_ (.A1(_01648_),
    .A2(_01687_),
    .A3(_01666_),
    .B1(_01745_),
    .C1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01746_));
 sky130_fd_sc_hd__nand2_1 _07066_ (.A(_01590_),
    .B(_01733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01747_));
 sky130_fd_sc_hd__or3_1 _07067_ (.A(_01649_),
    .B(_01602_),
    .C(_01694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01748_));
 sky130_fd_sc_hd__a21oi_1 _07068_ (.A1(_01747_),
    .A2(_01748_),
    .B1(_01644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01749_));
 sky130_fd_sc_hd__or2_1 _07069_ (.A(_00454_),
    .B(_01600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01750_));
 sky130_fd_sc_hd__a21oi_2 _07070_ (.A1(_01606_),
    .A2(_01750_),
    .B1(_01639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01751_));
 sky130_fd_sc_hd__o21a_1 _07071_ (.A1(_01595_),
    .A2(_01751_),
    .B1(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01752_));
 sky130_fd_sc_hd__a41o_1 _07072_ (.A1(_01625_),
    .A2(_01620_),
    .A3(_01653_),
    .A4(_01635_),
    .B1(_01752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01753_));
 sky130_fd_sc_hd__o21a_1 _07073_ (.A1(_01749_),
    .A2(_01753_),
    .B1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01754_));
 sky130_fd_sc_hd__a31o_1 _07074_ (.A1(_00457_),
    .A2(_01742_),
    .A3(_01746_),
    .B1(_01754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00030_));
 sky130_fd_sc_hd__a311o_1 _07075_ (.A1(_00455_),
    .A2(_01750_),
    .A3(_01680_),
    .B1(_01715_),
    .C1(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01755_));
 sky130_fd_sc_hd__a211o_1 _07076_ (.A1(_01648_),
    .A2(_01687_),
    .B1(_01628_),
    .C1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01756_));
 sky130_fd_sc_hd__or2_1 _07077_ (.A(_01632_),
    .B(_01615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01757_));
 sky130_fd_sc_hd__a21o_1 _07078_ (.A1(_01722_),
    .A2(_01757_),
    .B1(_01644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01758_));
 sky130_fd_sc_hd__or3_1 _07079_ (.A(_01632_),
    .B(_01617_),
    .C(_01721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01759_));
 sky130_fd_sc_hd__a21oi_1 _07080_ (.A1(_01758_),
    .A2(_01759_),
    .B1(_01631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01760_));
 sky130_fd_sc_hd__a31o_1 _07081_ (.A1(_00457_),
    .A2(_01755_),
    .A3(_01756_),
    .B1(_01760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00031_));
 sky130_fd_sc_hd__nor2_1 _07082_ (.A(_01602_),
    .B(_01609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_1 _07083_ (.A(_01643_),
    .B(_01602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01762_));
 sky130_fd_sc_hd__o21ai_1 _07084_ (.A1(_01694_),
    .A2(_01762_),
    .B1(_01620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01763_));
 sky130_fd_sc_hd__or2_1 _07085_ (.A(_01761_),
    .B(_01763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01764_));
 sky130_fd_sc_hd__a211o_1 _07086_ (.A1(_01721_),
    .A2(_01701_),
    .B1(_01621_),
    .C1(_01616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01765_));
 sky130_fd_sc_hd__nand2_1 _07087_ (.A(_01637_),
    .B(_01591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01766_));
 sky130_fd_sc_hd__a21o_1 _07088_ (.A1(_01766_),
    .A2(_01762_),
    .B1(_01617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01767_));
 sky130_fd_sc_hd__nor2_1 _07089_ (.A(_01657_),
    .B(_01611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01768_));
 sky130_fd_sc_hd__a211o_1 _07090_ (.A1(_01768_),
    .A2(_01761_),
    .B1(_01751_),
    .C1(_01620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01769_));
 sky130_fd_sc_hd__and3_1 _07091_ (.A(_01663_),
    .B(_01767_),
    .C(_01769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01770_));
 sky130_fd_sc_hd__a31o_1 _07092_ (.A1(_00457_),
    .A2(_01764_),
    .A3(_01765_),
    .B1(_01770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00001_));
 sky130_fd_sc_hd__a32o_1 _07093_ (.A1(_01690_),
    .A2(_01625_),
    .A3(_01603_),
    .B1(_01682_),
    .B2(_01654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01771_));
 sky130_fd_sc_hd__a21oi_1 _07094_ (.A1(_01605_),
    .A2(_01647_),
    .B1(_01650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01772_));
 sky130_fd_sc_hd__or3_1 _07095_ (.A(_01657_),
    .B(_01646_),
    .C(_01696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01773_));
 sky130_fd_sc_hd__a22o_1 _07096_ (.A1(_01618_),
    .A2(_01771_),
    .B1(_01772_),
    .B2(_01773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01774_));
 sky130_fd_sc_hd__nor2_1 _07097_ (.A(_01646_),
    .B(_01634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _07098_ (.A(_01578_),
    .B(_01653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01776_));
 sky130_fd_sc_hd__a211o_1 _07099_ (.A1(_01654_),
    .A2(_01653_),
    .B1(_01776_),
    .C1(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01777_));
 sky130_fd_sc_hd__o311a_1 _07100_ (.A1(_01595_),
    .A2(_01729_),
    .A3(_01775_),
    .B1(_01777_),
    .C1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01778_));
 sky130_fd_sc_hd__a21o_1 _07101_ (.A1(_01679_),
    .A2(_01774_),
    .B1(_01778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00002_));
 sky130_fd_sc_hd__a21oi_1 _07102_ (.A1(_01622_),
    .A2(_01647_),
    .B1(_01710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01779_));
 sky130_fd_sc_hd__and3_1 _07103_ (.A(_01648_),
    .B(_01639_),
    .C(_01634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01780_));
 sky130_fd_sc_hd__o31ai_1 _07104_ (.A1(_01622_),
    .A2(_01687_),
    .A3(_01694_),
    .B1(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01781_));
 sky130_fd_sc_hd__o32a_1 _07105_ (.A1(_01644_),
    .A2(_01688_),
    .A3(_01779_),
    .B1(_01780_),
    .B2(_01781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01782_));
 sky130_fd_sc_hd__nor2_1 _07106_ (.A(_01743_),
    .B(_01647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01783_));
 sky130_fd_sc_hd__a31o_1 _07107_ (.A1(_01603_),
    .A2(_01594_),
    .A3(_01666_),
    .B1(_01617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01784_));
 sky130_fd_sc_hd__a31o_1 _07108_ (.A1(_01657_),
    .A2(_01580_),
    .A3(_01653_),
    .B1(_01734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01785_));
 sky130_fd_sc_hd__o211a_1 _07109_ (.A1(_01783_),
    .A2(_01784_),
    .B1(_01629_),
    .C1(_01785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01786_));
 sky130_fd_sc_hd__a21o_1 _07110_ (.A1(_01679_),
    .A2(_01782_),
    .B1(_01786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00003_));
 sky130_fd_sc_hd__o21a_1 _07111_ (.A1(_01649_),
    .A2(_01696_),
    .B1(_01603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01787_));
 sky130_fd_sc_hd__a211o_1 _07112_ (.A1(_01682_),
    .A2(_01706_),
    .B1(_01787_),
    .C1(_01644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01788_));
 sky130_fd_sc_hd__a21o_1 _07113_ (.A1(_01701_),
    .A2(_01704_),
    .B1(_01705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01789_));
 sky130_fd_sc_hd__or2_1 _07114_ (.A(_01620_),
    .B(_01780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01790_));
 sky130_fd_sc_hd__a31o_1 _07115_ (.A1(_01578_),
    .A2(_01690_),
    .A3(_01703_),
    .B1(_01790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01791_));
 sky130_fd_sc_hd__nand2_1 _07116_ (.A(_01637_),
    .B(_01642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01792_));
 sky130_fd_sc_hd__o22a_1 _07117_ (.A1(_01792_),
    .A2(_01653_),
    .B1(_01626_),
    .B2(_01659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01793_));
 sky130_fd_sc_hd__a21oi_1 _07118_ (.A1(_00456_),
    .A2(_01793_),
    .B1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01794_));
 sky130_fd_sc_hd__a32o_1 _07119_ (.A1(_01631_),
    .A2(_01788_),
    .A3(_01789_),
    .B1(_01791_),
    .B2(_01794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00004_));
 sky130_fd_sc_hd__nand2_1 _07120_ (.A(_01617_),
    .B(_01727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_1 _07121_ (.A(_01640_),
    .B(_01594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _07122_ (.A(_01719_),
    .B(_01673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01797_));
 sky130_fd_sc_hd__or2_1 _07123_ (.A(_01584_),
    .B(_01797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01798_));
 sky130_fd_sc_hd__nor2_1 _07124_ (.A(_01657_),
    .B(_01627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01799_));
 sky130_fd_sc_hd__o32a_1 _07125_ (.A1(_01761_),
    .A2(_01795_),
    .A3(_01796_),
    .B1(_01798_),
    .B2(_01799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01800_));
 sky130_fd_sc_hd__o221a_1 _07126_ (.A1(_01719_),
    .A2(_01641_),
    .B1(_01696_),
    .B2(_01659_),
    .C1(_00456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01801_));
 sky130_fd_sc_hd__a31o_1 _07127_ (.A1(_01642_),
    .A2(_01647_),
    .A3(_01594_),
    .B1(_01726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01802_));
 sky130_fd_sc_hd__nand2_1 _07128_ (.A(_01631_),
    .B(_01802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01803_));
 sky130_fd_sc_hd__o22a_1 _07129_ (.A1(_01631_),
    .A2(_01800_),
    .B1(_01801_),
    .B2(_01803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00005_));
 sky130_fd_sc_hd__nor2_1 _07130_ (.A(_01632_),
    .B(_01659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01804_));
 sky130_fd_sc_hd__a311o_1 _07131_ (.A1(_01593_),
    .A2(_01648_),
    .A3(_01659_),
    .B1(_01804_),
    .C1(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01805_));
 sky130_fd_sc_hd__o31a_1 _07132_ (.A1(_01667_),
    .A2(_01583_),
    .A3(_01640_),
    .B1(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01806_));
 sky130_fd_sc_hd__o311a_1 _07133_ (.A1(_01632_),
    .A2(_01584_),
    .A3(_01673_),
    .B1(_01805_),
    .C1(_01806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01807_));
 sky130_fd_sc_hd__a21oi_1 _07134_ (.A1(_01666_),
    .A2(_01706_),
    .B1(_01646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01808_));
 sky130_fd_sc_hd__a21oi_1 _07135_ (.A1(_01578_),
    .A2(_01612_),
    .B1(_01640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01809_));
 sky130_fd_sc_hd__o221a_1 _07136_ (.A1(_01705_),
    .A2(_01808_),
    .B1(_01809_),
    .B2(_01598_),
    .C1(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01810_));
 sky130_fd_sc_hd__or2_1 _07137_ (.A(_01807_),
    .B(_01810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01811_));
 sky130_fd_sc_hd__clkbuf_1 _07138_ (.A(_01811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00006_));
 sky130_fd_sc_hd__and3_1 _07139_ (.A(_01585_),
    .B(_00455_),
    .C(_01681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01812_));
 sky130_fd_sc_hd__a311o_1 _07140_ (.A1(_01644_),
    .A2(_01610_),
    .A3(_01660_),
    .B1(_01797_),
    .C1(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01813_));
 sky130_fd_sc_hd__a21oi_1 _07141_ (.A1(_01594_),
    .A2(_01666_),
    .B1(_00455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01814_));
 sky130_fd_sc_hd__a221o_1 _07142_ (.A1(_01612_),
    .A2(_01703_),
    .B1(_01721_),
    .B2(_01719_),
    .C1(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01815_));
 sky130_fd_sc_hd__o21ai_1 _07143_ (.A1(_01705_),
    .A2(_01814_),
    .B1(_01815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01816_));
 sky130_fd_sc_hd__o22a_1 _07144_ (.A1(_01812_),
    .A2(_01813_),
    .B1(_01816_),
    .B2(_00457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00007_));
 sky130_fd_sc_hd__a21o_1 _07145_ (.A1(_00455_),
    .A2(_01739_),
    .B1(_01798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01817_));
 sky130_fd_sc_hd__a211o_1 _07146_ (.A1(_01710_),
    .A2(_01687_),
    .B1(_01714_),
    .C1(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01818_));
 sky130_fd_sc_hd__and3_1 _07147_ (.A(_01690_),
    .B(_01750_),
    .C(_01682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01819_));
 sky130_fd_sc_hd__and2_1 _07148_ (.A(_01743_),
    .B(_01639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01820_));
 sky130_fd_sc_hd__a311o_1 _07149_ (.A1(_01603_),
    .A2(_01610_),
    .A3(_01706_),
    .B1(_01820_),
    .C1(_01620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01821_));
 sky130_fd_sc_hd__o311a_1 _07150_ (.A1(_01650_),
    .A2(_01728_),
    .A3(_01819_),
    .B1(_01821_),
    .C1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01822_));
 sky130_fd_sc_hd__a31o_1 _07151_ (.A1(_01679_),
    .A2(_01817_),
    .A3(_01818_),
    .B1(_01822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00008_));
 sky130_fd_sc_hd__nor2_1 _07152_ (.A(_01652_),
    .B(_01819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01823_));
 sky130_fd_sc_hd__nand2_1 _07153_ (.A(_01667_),
    .B(_01640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01824_));
 sky130_fd_sc_hd__or3b_1 _07154_ (.A(_01601_),
    .B(_01658_),
    .C_N(_01824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01825_));
 sky130_fd_sc_hd__a32o_1 _07155_ (.A1(_00456_),
    .A2(_01610_),
    .A3(_01773_),
    .B1(_01823_),
    .B2(_01825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01826_));
 sky130_fd_sc_hd__a31o_1 _07156_ (.A1(_01578_),
    .A2(_01625_),
    .A3(_01703_),
    .B1(_01790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01827_));
 sky130_fd_sc_hd__a31o_1 _07157_ (.A1(_01607_),
    .A2(_01690_),
    .A3(_01766_),
    .B1(_01700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01828_));
 sky130_fd_sc_hd__o21a_1 _07158_ (.A1(_01618_),
    .A2(_01828_),
    .B1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01829_));
 sky130_fd_sc_hd__a2bb2o_1 _07159_ (.A1_N(_00457_),
    .A2_N(_01826_),
    .B1(_01827_),
    .B2(_01829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00009_));
 sky130_fd_sc_hd__nor2_1 _07160_ (.A(_00454_),
    .B(_00452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01830_));
 sky130_fd_sc_hd__a21o_1 _07161_ (.A1(_01639_),
    .A2(_01696_),
    .B1(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01831_));
 sky130_fd_sc_hd__o32a_1 _07162_ (.A1(_01583_),
    .A2(_01830_),
    .A3(_01674_),
    .B1(_01738_),
    .B2(_01831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01832_));
 sky130_fd_sc_hd__inv_1 _07163_ (.A(_01832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01833_));
 sky130_fd_sc_hd__o32a_1 _07164_ (.A1(_01580_),
    .A2(_01602_),
    .A3(_01830_),
    .B1(_01747_),
    .B2(_01608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01834_));
 sky130_fd_sc_hd__o22a_1 _07165_ (.A1(_01703_),
    .A2(_01831_),
    .B1(_01834_),
    .B2(_01617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _07166_ (.A0(_01833_),
    .A1(_01835_),
    .S(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01836_));
 sky130_fd_sc_hd__clkbuf_1 _07167_ (.A(_01836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00010_));
 sky130_fd_sc_hd__o31a_1 _07168_ (.A1(_01657_),
    .A2(_01646_),
    .A3(_01611_),
    .B1(_01661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01837_));
 sky130_fd_sc_hd__o22a_1 _07169_ (.A1(_01790_),
    .A2(_01796_),
    .B1(_01837_),
    .B2(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01838_));
 sky130_fd_sc_hd__o21ba_1 _07170_ (.A1(_01636_),
    .A2(_01682_),
    .B1_N(_01729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01839_));
 sky130_fd_sc_hd__nor2_1 _07171_ (.A(_01830_),
    .B(_01658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01840_));
 sky130_fd_sc_hd__o221a_1 _07172_ (.A1(_01694_),
    .A2(_01762_),
    .B1(_01840_),
    .B2(_01703_),
    .C1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01841_));
 sky130_fd_sc_hd__or3_1 _07173_ (.A(_01570_),
    .B(_01839_),
    .C(_01841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01842_));
 sky130_fd_sc_hd__o21ai_1 _07174_ (.A1(_01631_),
    .A2(_01838_),
    .B1(_01842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00012_));
 sky130_fd_sc_hd__a211o_1 _07175_ (.A1(_01591_),
    .A2(_01666_),
    .B1(_01787_),
    .C1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01843_));
 sky130_fd_sc_hd__o32a_1 _07176_ (.A1(_01608_),
    .A2(_01581_),
    .A3(_01626_),
    .B1(_01653_),
    .B2(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01844_));
 sky130_fd_sc_hd__or2_1 _07177_ (.A(_01621_),
    .B(_01844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01845_));
 sky130_fd_sc_hd__a211o_1 _07178_ (.A1(_01591_),
    .A2(_01612_),
    .B1(_01776_),
    .C1(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01846_));
 sky130_fd_sc_hd__o311a_1 _07179_ (.A1(_01650_),
    .A2(_01714_),
    .A3(_01820_),
    .B1(_01846_),
    .C1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01847_));
 sky130_fd_sc_hd__a31o_1 _07180_ (.A1(_00457_),
    .A2(_01843_),
    .A3(_01845_),
    .B1(_01847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00013_));
 sky130_fd_sc_hd__a221o_1 _07181_ (.A1(_01687_),
    .A2(_01719_),
    .B1(_01702_),
    .B2(_01703_),
    .C1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01848_));
 sky130_fd_sc_hd__nand2_1 _07182_ (.A(_00452_),
    .B(_01640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01849_));
 sky130_fd_sc_hd__a221o_1 _07183_ (.A1(_01657_),
    .A2(_01687_),
    .B1(_01849_),
    .B2(_01633_),
    .C1(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01850_));
 sky130_fd_sc_hd__a21oi_1 _07184_ (.A1(_01792_),
    .A2(_01634_),
    .B1(_01653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01851_));
 sky130_fd_sc_hd__a311o_1 _07185_ (.A1(_01637_),
    .A2(_01603_),
    .A3(_01701_),
    .B1(_01775_),
    .C1(_01620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01852_));
 sky130_fd_sc_hd__o311a_1 _07186_ (.A1(_01650_),
    .A2(_01681_),
    .A3(_01851_),
    .B1(_01852_),
    .C1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01853_));
 sky130_fd_sc_hd__a31o_1 _07187_ (.A1(_01679_),
    .A2(_01848_),
    .A3(_01850_),
    .B1(_01853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00014_));
 sky130_fd_sc_hd__or3b_1 _07188_ (.A(_01808_),
    .B(_01650_),
    .C_N(_01627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01854_));
 sky130_fd_sc_hd__a21o_1 _07189_ (.A1(_01792_),
    .A2(_01703_),
    .B1(_01598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01855_));
 sky130_fd_sc_hd__o22a_1 _07190_ (.A1(_01622_),
    .A2(_01696_),
    .B1(_01747_),
    .B2(_01611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01856_));
 sky130_fd_sc_hd__a311o_1 _07191_ (.A1(_01665_),
    .A2(_01647_),
    .A3(_01626_),
    .B1(_01856_),
    .C1(_01650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01857_));
 sky130_fd_sc_hd__a31oi_1 _07192_ (.A1(_01618_),
    .A2(_01748_),
    .A3(_01744_),
    .B1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01858_));
 sky130_fd_sc_hd__a32o_1 _07193_ (.A1(_01631_),
    .A2(_01854_),
    .A3(_01855_),
    .B1(_01857_),
    .B2(_01858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00015_));
 sky130_fd_sc_hd__o21ai_1 _07194_ (.A1(_01622_),
    .A2(_01603_),
    .B1(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01859_));
 sky130_fd_sc_hd__a31o_1 _07195_ (.A1(_01647_),
    .A2(_01610_),
    .A3(_01706_),
    .B1(_01859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01860_));
 sky130_fd_sc_hd__a31o_1 _07196_ (.A1(_01665_),
    .A2(_01647_),
    .A3(_01733_),
    .B1(_01598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01861_));
 sky130_fd_sc_hd__a21oi_1 _07197_ (.A1(_01623_),
    .A2(_01723_),
    .B1(_01611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01862_));
 sky130_fd_sc_hd__or3_1 _07198_ (.A(_01584_),
    .B(_01849_),
    .C(_01658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01863_));
 sky130_fd_sc_hd__o211a_1 _07199_ (.A1(_01644_),
    .A2(_01862_),
    .B1(_01863_),
    .C1(_01571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01864_));
 sky130_fd_sc_hd__a31oi_1 _07200_ (.A1(_01679_),
    .A2(_01860_),
    .A3(_01861_),
    .B1(_01864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00016_));
 sky130_fd_sc_hd__a211o_1 _07201_ (.A1(_00455_),
    .A2(_01696_),
    .B1(_01689_),
    .C1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01865_));
 sky130_fd_sc_hd__a211o_1 _07202_ (.A1(_01600_),
    .A2(_01682_),
    .B1(_01694_),
    .C1(_01649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01866_));
 sky130_fd_sc_hd__nand2_1 _07203_ (.A(_01823_),
    .B(_01866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01867_));
 sky130_fd_sc_hd__and3_1 _07204_ (.A(_01593_),
    .B(_01646_),
    .C(_01750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01868_));
 sky130_fd_sc_hd__o21ai_1 _07205_ (.A1(_01804_),
    .A2(_01868_),
    .B1(_01644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01869_));
 sky130_fd_sc_hd__o211a_1 _07206_ (.A1(_01745_),
    .A2(_01831_),
    .B1(_01869_),
    .C1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01870_));
 sky130_fd_sc_hd__a31o_1 _07207_ (.A1(_00457_),
    .A2(_01865_),
    .A3(_01867_),
    .B1(_01870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00017_));
 sky130_fd_sc_hd__a21oi_1 _07208_ (.A1(_01643_),
    .A2(_01610_),
    .B1(_01647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _07209_ (.A(_01608_),
    .B(_01602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01872_));
 sky130_fd_sc_hd__o31a_1 _07210_ (.A1(_01622_),
    .A2(_01639_),
    .A3(_01658_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01873_));
 sky130_fd_sc_hd__a21bo_1 _07211_ (.A1(_01593_),
    .A2(_01872_),
    .B1_N(_01873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01874_));
 sky130_fd_sc_hd__o31a_1 _07212_ (.A1(_01650_),
    .A2(_01851_),
    .A3(_01871_),
    .B1(_01874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01875_));
 sky130_fd_sc_hd__o21a_1 _07213_ (.A1(_01581_),
    .A2(_01655_),
    .B1(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01876_));
 sky130_fd_sc_hd__a31o_1 _07214_ (.A1(_01690_),
    .A2(_01687_),
    .A3(_01609_),
    .B1(_01685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01877_));
 sky130_fd_sc_hd__o21ai_1 _07215_ (.A1(_01618_),
    .A2(_01877_),
    .B1(_01679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01878_));
 sky130_fd_sc_hd__o22a_1 _07216_ (.A1(_01679_),
    .A2(_01875_),
    .B1(_01876_),
    .B2(_01878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00018_));
 sky130_fd_sc_hd__o31ai_1 _07217_ (.A1(_01595_),
    .A2(_01604_),
    .A3(_01751_),
    .B1(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01879_));
 sky130_fd_sc_hd__a211o_1 _07218_ (.A1(_01684_),
    .A2(_01820_),
    .B1(_01799_),
    .C1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01880_));
 sky130_fd_sc_hd__o2bb2a_1 _07219_ (.A1_N(_01733_),
    .A2_N(_01659_),
    .B1(_01690_),
    .B2(_01603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01881_));
 sky130_fd_sc_hd__or3_1 _07220_ (.A(_01584_),
    .B(_01796_),
    .C(_01872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01882_));
 sky130_fd_sc_hd__o211a_1 _07221_ (.A1(_00456_),
    .A2(_01881_),
    .B1(_01882_),
    .C1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01883_));
 sky130_fd_sc_hd__a31o_1 _07222_ (.A1(_01631_),
    .A2(_01879_),
    .A3(_01880_),
    .B1(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00019_));
 sky130_fd_sc_hd__a21oi_1 _07223_ (.A1(_01593_),
    .A2(_01648_),
    .B1(_01647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01884_));
 sky130_fd_sc_hd__or3_1 _07224_ (.A(_01650_),
    .B(_01745_),
    .C(_01884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01885_));
 sky130_fd_sc_hd__a221o_1 _07225_ (.A1(_01643_),
    .A2(_00455_),
    .B1(_01604_),
    .B2(_01701_),
    .C1(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01886_));
 sky130_fd_sc_hd__or3_1 _07226_ (.A(_01620_),
    .B(_01628_),
    .C(_01872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01887_));
 sky130_fd_sc_hd__o311a_1 _07227_ (.A1(_01650_),
    .A2(_01700_),
    .A3(_01711_),
    .B1(_01887_),
    .C1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01888_));
 sky130_fd_sc_hd__a31o_1 _07228_ (.A1(_01631_),
    .A2(_01885_),
    .A3(_01886_),
    .B1(_01888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00020_));
 sky130_fd_sc_hd__o211a_1 _07229_ (.A1(_01632_),
    .A2(_01615_),
    .B1(_01673_),
    .C1(_01618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01889_));
 sky130_fd_sc_hd__o21ai_1 _07230_ (.A1(_00454_),
    .A2(_01637_),
    .B1(_01682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01890_));
 sky130_fd_sc_hd__a31o_1 _07231_ (.A1(_01621_),
    .A2(_01615_),
    .A3(_01890_),
    .B1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01891_));
 sky130_fd_sc_hd__and3_1 _07232_ (.A(_01665_),
    .B(_01648_),
    .C(_01809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01892_));
 sky130_fd_sc_hd__o21ai_1 _07233_ (.A1(_01739_),
    .A2(_01809_),
    .B1(_00456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01893_));
 sky130_fd_sc_hd__o211a_1 _07234_ (.A1(_01607_),
    .A2(_01580_),
    .B1(_01646_),
    .C1(_00452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01894_));
 sky130_fd_sc_hd__o31a_1 _07235_ (.A1(_01652_),
    .A2(_01761_),
    .A3(_01894_),
    .B1(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01895_));
 sky130_fd_sc_hd__o21ai_1 _07236_ (.A1(_01892_),
    .A2(_01893_),
    .B1(_01895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01896_));
 sky130_fd_sc_hd__o21ai_1 _07237_ (.A1(_01889_),
    .A2(_01891_),
    .B1(_01896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00021_));
 sky130_fd_sc_hd__a211o_1 _07238_ (.A1(_01849_),
    .A2(_01633_),
    .B1(_01611_),
    .C1(_01657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01897_));
 sky130_fd_sc_hd__or2_1 _07239_ (.A(_01724_),
    .B(_01897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01898_));
 sky130_fd_sc_hd__nand2_1 _07240_ (.A(_01724_),
    .B(_01897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01899_));
 sky130_fd_sc_hd__a31o_1 _07241_ (.A1(_01653_),
    .A2(_01768_),
    .A3(_01684_),
    .B1(_01763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01900_));
 sky130_fd_sc_hd__o211a_1 _07242_ (.A1(_01668_),
    .A2(_01795_),
    .B1(_01900_),
    .C1(_01663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01901_));
 sky130_fd_sc_hd__a31o_1 _07243_ (.A1(_01631_),
    .A2(_01898_),
    .A3(_01899_),
    .B1(_01901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00023_));
 sky130_fd_sc_hd__a21o_1 _07244_ (.A1(_00455_),
    .A2(_01680_),
    .B1(_01798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01902_));
 sky130_fd_sc_hd__a211o_1 _07245_ (.A1(_00454_),
    .A2(_01824_),
    .B1(_01783_),
    .C1(_01621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01903_));
 sky130_fd_sc_hd__a21oi_1 _07246_ (.A1(_01613_),
    .A2(_01695_),
    .B1(_01644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01904_));
 sky130_fd_sc_hd__o21a_1 _07247_ (.A1(_01752_),
    .A2(_01904_),
    .B1(_01629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01905_));
 sky130_fd_sc_hd__a31o_1 _07248_ (.A1(_01679_),
    .A2(_01902_),
    .A3(_01903_),
    .B1(_01905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00024_));
 sky130_fd_sc_hd__or3_1 _07249_ (.A(\state[2] ),
    .B(_00032_),
    .C(_01563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01906_));
 sky130_fd_sc_hd__and2_1 _07250_ (.A(\sha256cu.byte_stop ),
    .B(_01906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01907_));
 sky130_fd_sc_hd__clkbuf_1 _07251_ (.A(_01907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00068_));
 sky130_fd_sc_hd__a31o_1 _07252_ (.A1(\state[1] ),
    .A2(\sha256cu.hashing_done ),
    .A3(_01560_),
    .B1(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01908_));
 sky130_fd_sc_hd__and2b_1 _07253_ (.A_N(net257),
    .B(_01908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01909_));
 sky130_fd_sc_hd__clkbuf_1 _07254_ (.A(_01909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00069_));
 sky130_fd_sc_hd__o21ba_1 _07255_ (.A1(net259),
    .A2(\state[3] ),
    .B1_N(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00070_));
 sky130_fd_sc_hd__inv_2 _07256_ (.A(\state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01910_));
 sky130_fd_sc_hd__clkinv_4 _07257_ (.A(_01564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01911_));
 sky130_fd_sc_hd__buf_4 _07258_ (.A(_01911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01912_));
 sky130_fd_sc_hd__buf_6 _07259_ (.A(_01912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01913_));
 sky130_fd_sc_hd__a311oi_1 _07260_ (.A1(\state[1] ),
    .A2(\sha256cu.hashing_done ),
    .A3(_01910_),
    .B1(net257),
    .C1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00071_));
 sky130_fd_sc_hd__and2_1 _07261_ (.A(\sha256cu.m_pad_pars.add_512_block[5] ),
    .B(\sha256cu.m_pad_pars.add_512_block[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01914_));
 sky130_fd_sc_hd__a31o_1 _07262_ (.A1(\sha256cu.m_pad_pars.add_512_block[2] ),
    .A2(\sha256cu.m_pad_pars.add_512_block[1] ),
    .A3(\sha256cu.m_pad_pars.add_512_block[0] ),
    .B1(\sha256cu.m_pad_pars.add_512_block[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01915_));
 sky130_fd_sc_hd__a21oi_2 _07263_ (.A1(_01914_),
    .A2(_01915_),
    .B1(\sha256cu.m_pad_pars.add_512_block[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01916_));
 sky130_fd_sc_hd__or2b_1 _07264_ (.A(\sha256cu.byte_rdy ),
    .B_N(\sha256cu.byte_stop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01917_));
 sky130_fd_sc_hd__or2_1 _07265_ (.A(_01916_),
    .B(_01917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01918_));
 sky130_fd_sc_hd__clkbuf_4 _07266_ (.A(_01918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01919_));
 sky130_fd_sc_hd__buf_4 _07267_ (.A(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01920_));
 sky130_fd_sc_hd__clkbuf_4 _07268_ (.A(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01921_));
 sky130_fd_sc_hd__or2_1 _07269_ (.A(_01911_),
    .B(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01922_));
 sky130_fd_sc_hd__clkbuf_4 _07270_ (.A(_01922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01923_));
 sky130_fd_sc_hd__clkbuf_2 _07271_ (.A(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01924_));
 sky130_fd_sc_hd__and2_1 _07272_ (.A(\sha256cu.m_pad_pars.block_512[63][0] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01925_));
 sky130_fd_sc_hd__clkbuf_1 _07273_ (.A(_01925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00072_));
 sky130_fd_sc_hd__and2_1 _07274_ (.A(\sha256cu.m_pad_pars.block_512[63][1] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01926_));
 sky130_fd_sc_hd__clkbuf_1 _07275_ (.A(_01926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00073_));
 sky130_fd_sc_hd__and2_1 _07276_ (.A(\sha256cu.m_pad_pars.block_512[63][2] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01927_));
 sky130_fd_sc_hd__clkbuf_1 _07277_ (.A(_01927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00074_));
 sky130_fd_sc_hd__clkbuf_4 _07278_ (.A(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _07279_ (.A0(\sha256cu.m_pad_pars.m_size[3] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][3] ),
    .S(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01929_));
 sky130_fd_sc_hd__clkbuf_1 _07280_ (.A(_01929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _07281_ (.A0(\sha256cu.m_pad_pars.m_size[4] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][4] ),
    .S(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01930_));
 sky130_fd_sc_hd__clkbuf_1 _07282_ (.A(_01930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _07283_ (.A0(\sha256cu.m_pad_pars.m_size[5] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][5] ),
    .S(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01931_));
 sky130_fd_sc_hd__clkbuf_1 _07284_ (.A(_01931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _07285_ (.A0(\sha256cu.m_pad_pars.m_size[6] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][6] ),
    .S(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01932_));
 sky130_fd_sc_hd__clkbuf_1 _07286_ (.A(_01932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _07287_ (.A0(\sha256cu.m_pad_pars.m_size[7] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][7] ),
    .S(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01933_));
 sky130_fd_sc_hd__clkbuf_1 _07288_ (.A(_01933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00079_));
 sky130_fd_sc_hd__or2b_1 _07289_ (.A(\sha256cu.byte_rdy ),
    .B_N(_01906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01934_));
 sky130_fd_sc_hd__clkbuf_1 _07290_ (.A(_01934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00080_));
 sky130_fd_sc_hd__nor2_2 _07291_ (.A(\sha256cu.m_pad_pars.add_out0[3] ),
    .B(\sha256cu.m_pad_pars.add_out0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_2 _07292_ (.A(\sha256cu.m_pad_pars.add_out0[5] ),
    .B(\sha256cu.m_pad_pars.add_out0[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_2 _07293_ (.A(_01935_),
    .B(_01936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01937_));
 sky130_fd_sc_hd__o21a_1 _07294_ (.A1(\sha256cu.m_pad_pars.add_out0[6] ),
    .A2(_01937_),
    .B1(\sha256cu.m_pad_pars.add_out3[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01938_));
 sky130_fd_sc_hd__clkbuf_4 _07295_ (.A(\sha256cu.m_pad_pars.add_512_block[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01939_));
 sky130_fd_sc_hd__or2_2 _07296_ (.A(\sha256cu.m_pad_pars.add_512_block[3] ),
    .B(\sha256cu.m_pad_pars.add_512_block[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01940_));
 sky130_fd_sc_hd__or2_2 _07297_ (.A(\sha256cu.m_pad_pars.add_512_block[1] ),
    .B(_01939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01941_));
 sky130_fd_sc_hd__nor2_4 _07298_ (.A(_01940_),
    .B(_01941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01942_));
 sky130_fd_sc_hd__or2_2 _07299_ (.A(\sha256cu.m_pad_pars.add_512_block[5] ),
    .B(\sha256cu.m_pad_pars.add_512_block[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01943_));
 sky130_fd_sc_hd__clkinv_2 _07300_ (.A(_01943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_2 _07301_ (.A(\sha256cu.byte_stop ),
    .B(_01916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01945_));
 sky130_fd_sc_hd__a21oi_1 _07302_ (.A1(_01942_),
    .A2(_01944_),
    .B1(_01945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01946_));
 sky130_fd_sc_hd__a21o_1 _07303_ (.A1(\sha256cu.byte_stop ),
    .A2(_01916_),
    .B1(\sha256cu.byte_rdy ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01947_));
 sky130_fd_sc_hd__nand2_1 _07304_ (.A(_01939_),
    .B(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01948_));
 sky130_fd_sc_hd__o31a_1 _07305_ (.A1(_01939_),
    .A2(\sha256cu.byte_rdy ),
    .A3(_01946_),
    .B1(_01948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01949_));
 sky130_fd_sc_hd__nand2_2 _07306_ (.A(\sha256cu.m_pad_pars.add_512_block[5] ),
    .B(\sha256cu.m_pad_pars.add_512_block[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01950_));
 sky130_fd_sc_hd__or2_1 _07307_ (.A(\sha256cu.m_pad_pars.add_512_block[6] ),
    .B(_01950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01951_));
 sky130_fd_sc_hd__clkbuf_4 _07308_ (.A(_01951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01952_));
 sky130_fd_sc_hd__nand2b_2 _07309_ (.A_N(\sha256cu.m_pad_pars.add_512_block[3] ),
    .B(\sha256cu.m_pad_pars.add_512_block[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01953_));
 sky130_fd_sc_hd__or4b_1 _07310_ (.A(\sha256cu.byte_stop ),
    .B(_01952_),
    .C(_01953_),
    .D_N(\sha256cu.m_pad_pars.add_512_block[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01954_));
 sky130_fd_sc_hd__inv_2 _07311_ (.A(_01954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01955_));
 sky130_fd_sc_hd__clkinv_2 _07312_ (.A(\sha256cu.m_pad_pars.temp_chk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01956_));
 sky130_fd_sc_hd__a21oi_1 _07313_ (.A1(_01942_),
    .A2(_01944_),
    .B1(_01956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01957_));
 sky130_fd_sc_hd__o21ai_1 _07314_ (.A1(_01917_),
    .A2(_01957_),
    .B1(\sha256cu.iter_processing.padding_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01958_));
 sky130_fd_sc_hd__and2_1 _07315_ (.A(_01919_),
    .B(_01958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01959_));
 sky130_fd_sc_hd__a21o_1 _07316_ (.A1(_01949_),
    .A2(_01955_),
    .B1(_01959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01960_));
 sky130_fd_sc_hd__nor2_4 _07317_ (.A(_01938_),
    .B(_01960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01961_));
 sky130_fd_sc_hd__and2_1 _07318_ (.A(\sha256cu.m_pad_pars.add_out1[2] ),
    .B(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01962_));
 sky130_fd_sc_hd__clkbuf_4 _07319_ (.A(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01963_));
 sky130_fd_sc_hd__clkbuf_4 _07320_ (.A(_01564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01964_));
 sky130_fd_sc_hd__buf_6 _07321_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01965_));
 sky130_fd_sc_hd__buf_4 _07322_ (.A(_01965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01966_));
 sky130_fd_sc_hd__o21ai_1 _07323_ (.A1(\sha256cu.m_pad_pars.add_out1[2] ),
    .A2(_01963_),
    .B1(_01966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _07324_ (.A(_01962_),
    .B(_01967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _07325_ (.A(\sha256cu.m_pad_pars.add_out1[3] ),
    .B(\sha256cu.m_pad_pars.add_out1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01968_));
 sky130_fd_sc_hd__or2_2 _07326_ (.A(_01938_),
    .B(_01960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01969_));
 sky130_fd_sc_hd__clkbuf_8 _07327_ (.A(_01969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01970_));
 sky130_fd_sc_hd__buf_4 _07328_ (.A(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01971_));
 sky130_fd_sc_hd__buf_8 _07329_ (.A(_01564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01972_));
 sky130_fd_sc_hd__buf_4 _07330_ (.A(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01973_));
 sky130_fd_sc_hd__clkbuf_8 _07331_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01974_));
 sky130_fd_sc_hd__o221a_1 _07332_ (.A1(\sha256cu.m_pad_pars.add_out1[3] ),
    .A2(_01962_),
    .B1(_01968_),
    .B2(_01971_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00082_));
 sky130_fd_sc_hd__clkbuf_4 _07333_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01975_));
 sky130_fd_sc_hd__nand2_4 _07334_ (.A(_01564_),
    .B(_01969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01976_));
 sky130_fd_sc_hd__and2_2 _07335_ (.A(\sha256cu.m_pad_pars.add_out1[3] ),
    .B(\sha256cu.m_pad_pars.add_out1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01977_));
 sky130_fd_sc_hd__a21o_1 _07336_ (.A1(_01976_),
    .A2(_01977_),
    .B1(\sha256cu.m_pad_pars.add_out1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01978_));
 sky130_fd_sc_hd__nor2_1 _07337_ (.A(_01911_),
    .B(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01979_));
 sky130_fd_sc_hd__clkbuf_4 _07338_ (.A(_01979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01980_));
 sky130_fd_sc_hd__or3b_1 _07339_ (.A(_01980_),
    .B(_01968_),
    .C_N(\sha256cu.m_pad_pars.add_out1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01981_));
 sky130_fd_sc_hd__and3_1 _07340_ (.A(_01975_),
    .B(_01978_),
    .C(_01981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01982_));
 sky130_fd_sc_hd__clkbuf_1 _07341_ (.A(_01982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00083_));
 sky130_fd_sc_hd__buf_4 _07342_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01983_));
 sky130_fd_sc_hd__buf_4 _07343_ (.A(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01984_));
 sky130_fd_sc_hd__nor2b_2 _07344_ (.A(\sha256cu.m_pad_pars.add_out1[5] ),
    .B_N(\sha256cu.m_pad_pars.add_out1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01985_));
 sky130_fd_sc_hd__buf_4 _07345_ (.A(_01911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01986_));
 sky130_fd_sc_hd__nor2_4 _07346_ (.A(_01986_),
    .B(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01987_));
 sky130_fd_sc_hd__and3_1 _07347_ (.A(_01977_),
    .B(_01985_),
    .C(_01987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01988_));
 sky130_fd_sc_hd__a31o_1 _07348_ (.A1(\sha256cu.m_pad_pars.add_out1[5] ),
    .A2(_01984_),
    .A3(_01981_),
    .B1(_01988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00084_));
 sky130_fd_sc_hd__and2_1 _07349_ (.A(\sha256cu.m_pad_pars.add_out0[2] ),
    .B(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01989_));
 sky130_fd_sc_hd__o21ai_1 _07350_ (.A1(\sha256cu.m_pad_pars.add_out0[2] ),
    .A2(_01963_),
    .B1(_01966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_1 _07351_ (.A(_01989_),
    .B(_01990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00085_));
 sky130_fd_sc_hd__nand2_1 _07352_ (.A(\sha256cu.m_pad_pars.add_out0[3] ),
    .B(\sha256cu.m_pad_pars.add_out0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01991_));
 sky130_fd_sc_hd__o221a_1 _07353_ (.A1(\sha256cu.m_pad_pars.add_out0[3] ),
    .A2(_01989_),
    .B1(_01991_),
    .B2(_01971_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00086_));
 sky130_fd_sc_hd__and2_2 _07354_ (.A(\sha256cu.m_pad_pars.add_out0[3] ),
    .B(\sha256cu.m_pad_pars.add_out0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01992_));
 sky130_fd_sc_hd__and3_1 _07355_ (.A(\sha256cu.m_pad_pars.add_out0[4] ),
    .B(_01976_),
    .C(_01992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01993_));
 sky130_fd_sc_hd__buf_4 _07356_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01994_));
 sky130_fd_sc_hd__a21o_1 _07357_ (.A1(_01976_),
    .A2(_01992_),
    .B1(\sha256cu.m_pad_pars.add_out0[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01995_));
 sky130_fd_sc_hd__and3b_1 _07358_ (.A_N(_01993_),
    .B(_01994_),
    .C(_01995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01996_));
 sky130_fd_sc_hd__clkbuf_1 _07359_ (.A(_01996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00087_));
 sky130_fd_sc_hd__and3_1 _07360_ (.A(\sha256cu.m_pad_pars.add_out0[5] ),
    .B(\sha256cu.m_pad_pars.add_out0[4] ),
    .C(_01992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01997_));
 sky130_fd_sc_hd__clkbuf_4 _07361_ (.A(_01997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01998_));
 sky130_fd_sc_hd__nand2_1 _07362_ (.A(_01976_),
    .B(_01998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01999_));
 sky130_fd_sc_hd__buf_6 _07363_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02000_));
 sky130_fd_sc_hd__o211a_1 _07364_ (.A1(\sha256cu.m_pad_pars.add_out0[5] ),
    .A2(_01993_),
    .B1(_01999_),
    .C1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00088_));
 sky130_fd_sc_hd__and2_1 _07365_ (.A(_01976_),
    .B(_01998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02001_));
 sky130_fd_sc_hd__buf_4 _07366_ (.A(_01986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02002_));
 sky130_fd_sc_hd__a31o_1 _07367_ (.A1(\sha256cu.m_pad_pars.add_out0[6] ),
    .A2(_01963_),
    .A3(_01998_),
    .B1(_02002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02003_));
 sky130_fd_sc_hd__o21ba_1 _07368_ (.A1(\sha256cu.m_pad_pars.add_out0[6] ),
    .A2(_02001_),
    .B1_N(_02003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00089_));
 sky130_fd_sc_hd__or3b_1 _07369_ (.A(\sha256cu.counter_iteration[5] ),
    .B(\sha256cu.counter_iteration[4] ),
    .C_N(\sha256cu.counter_iteration[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02004_));
 sky130_fd_sc_hd__nor4_4 _07370_ (.A(\sha256cu.counter_iteration[3] ),
    .B(\sha256cu.counter_iteration[2] ),
    .C(\sha256cu.counter_iteration[1] ),
    .D(_02004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _07371_ (.A(\sha256cu.counter_iteration[0] ),
    .B(_02005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02006_));
 sky130_fd_sc_hd__and2_1 _07372_ (.A(_01964_),
    .B(\sha256cu.iter_processing.padding_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02007_));
 sky130_fd_sc_hd__a31o_1 _07373_ (.A1(\sha256cu.iter_processing.temp_case ),
    .A2(_02006_),
    .A3(_02007_),
    .B1(\sha256cu.iter_processing.temp_if ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00090_));
 sky130_fd_sc_hd__or4_1 _07374_ (.A(\sha256cu.counter_iteration[3] ),
    .B(\sha256cu.counter_iteration[2] ),
    .C(\sha256cu.counter_iteration[1] ),
    .D(_02004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02008_));
 sky130_fd_sc_hd__nor2_1 _07375_ (.A(\sha256cu.counter_iteration[0] ),
    .B(_02008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02009_));
 sky130_fd_sc_hd__and2b_1 _07376_ (.A_N(\sha256cu.m_out_digest.temp_delay ),
    .B(_02009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02010_));
 sky130_fd_sc_hd__xor2_1 _07377_ (.A(\sha256cu.m_out_digest.h_in[0] ),
    .B(\sha256cu.m_out_digest.H7[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02011_));
 sky130_fd_sc_hd__or4_1 _07378_ (.A(\sha256cu.counter_iteration[0] ),
    .B(\sha256cu.m_out_digest.temp_delay ),
    .C(_02008_),
    .D(_02011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02012_));
 sky130_fd_sc_hd__o211a_1 _07379_ (.A1(Hash_Digest),
    .A2(_02010_),
    .B1(_02012_),
    .C1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00091_));
 sky130_fd_sc_hd__o21a_1 _07380_ (.A1(\sha256cu.m_out_digest.temp_delay ),
    .A2(_02009_),
    .B1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _07381_ (.A0(\sha256cu.m_out_digest.H7[0] ),
    .A1(_02011_),
    .S(_02009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02013_));
 sky130_fd_sc_hd__or2_1 _07382_ (.A(_01913_),
    .B(_02013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02014_));
 sky130_fd_sc_hd__clkbuf_1 _07383_ (.A(_02014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00093_));
 sky130_fd_sc_hd__a22o_1 _07384_ (.A1(\sha256cu.iter_processing.temp_case ),
    .A2(_01984_),
    .B1(_02006_),
    .B2(_02007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00094_));
 sky130_fd_sc_hd__a21oi_2 _07385_ (.A1(\sha256cu.iter_processing.temp_case ),
    .A2(\sha256cu.iter_processing.padding_done ),
    .B1(\sha256cu.iter_processing.temp_if ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02015_));
 sky130_fd_sc_hd__or2_2 _07386_ (.A(_02005_),
    .B(_02015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02016_));
 sky130_fd_sc_hd__nand2_4 _07387_ (.A(_01564_),
    .B(_02016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02017_));
 sky130_fd_sc_hd__a21o_1 _07388_ (.A1(\sha256cu.m_out_digest.b_in[0] ),
    .A2(\sha256cu.m_out_digest.a_in[0] ),
    .B1(\sha256cu.m_out_digest.c_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02018_));
 sky130_fd_sc_hd__o21ai_1 _07389_ (.A1(\sha256cu.m_out_digest.b_in[0] ),
    .A2(\sha256cu.m_out_digest.a_in[0] ),
    .B1(_02018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02019_));
 sky130_fd_sc_hd__mux2_1 _07390_ (.A0(\sha256cu.m_out_digest.g_in[0] ),
    .A1(\sha256cu.m_out_digest.f_in[0] ),
    .S(\sha256cu.m_out_digest.e_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02020_));
 sky130_fd_sc_hd__xnor2_1 _07391_ (.A(_02019_),
    .B(_02020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02021_));
 sky130_fd_sc_hd__xnor2_1 _07392_ (.A(\sha256cu.iter_processing.w[0] ),
    .B(_02021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02022_));
 sky130_fd_sc_hd__xnor2_1 _07393_ (.A(\sha256cu.m_out_digest.e_in[11] ),
    .B(\sha256cu.m_out_digest.e_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02023_));
 sky130_fd_sc_hd__xnor2_2 _07394_ (.A(\sha256cu.m_out_digest.e_in[25] ),
    .B(_02023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02024_));
 sky130_fd_sc_hd__inv_2 _07395_ (.A(_02024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02025_));
 sky130_fd_sc_hd__buf_4 _07396_ (.A(\sha256cu.m_out_digest.a_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02026_));
 sky130_fd_sc_hd__clkbuf_4 _07397_ (.A(\sha256cu.m_out_digest.a_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02027_));
 sky130_fd_sc_hd__xnor2_1 _07398_ (.A(_02027_),
    .B(\sha256cu.m_out_digest.a_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02028_));
 sky130_fd_sc_hd__xnor2_2 _07399_ (.A(_02026_),
    .B(_02028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02029_));
 sky130_fd_sc_hd__xnor2_1 _07400_ (.A(\sha256cu.m_out_digest.h_in[0] ),
    .B(_02029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02030_));
 sky130_fd_sc_hd__xnor2_1 _07401_ (.A(_02025_),
    .B(_02030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02031_));
 sky130_fd_sc_hd__nor2_1 _07402_ (.A(_02022_),
    .B(_02031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02032_));
 sky130_fd_sc_hd__and2_1 _07403_ (.A(_02022_),
    .B(_02031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02033_));
 sky130_fd_sc_hd__nor2_1 _07404_ (.A(_02032_),
    .B(_02033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _07405_ (.A(\sha256cu.K[0] ),
    .B(_02034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02035_));
 sky130_fd_sc_hd__or2_1 _07406_ (.A(\sha256cu.K[0] ),
    .B(_02034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02036_));
 sky130_fd_sc_hd__buf_4 _07407_ (.A(_02016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02037_));
 sky130_fd_sc_hd__a32o_1 _07408_ (.A1(_02017_),
    .A2(_02035_),
    .A3(_02036_),
    .B1(_02037_),
    .B2(\sha256cu.m_out_digest.a_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02038_));
 sky130_fd_sc_hd__or2_1 _07409_ (.A(_01913_),
    .B(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02039_));
 sky130_fd_sc_hd__clkbuf_1 _07410_ (.A(_02039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00095_));
 sky130_fd_sc_hd__buf_4 _07411_ (.A(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02040_));
 sky130_fd_sc_hd__and2b_1 _07412_ (.A_N(_02019_),
    .B(_02020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02041_));
 sky130_fd_sc_hd__a21o_1 _07413_ (.A1(\sha256cu.iter_processing.w[0] ),
    .A2(_02021_),
    .B1(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02042_));
 sky130_fd_sc_hd__or2_1 _07414_ (.A(\sha256cu.m_out_digest.b_in[1] ),
    .B(\sha256cu.m_out_digest.a_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02043_));
 sky130_fd_sc_hd__a21o_1 _07415_ (.A1(\sha256cu.m_out_digest.b_in[1] ),
    .A2(\sha256cu.m_out_digest.a_in[1] ),
    .B1(\sha256cu.m_out_digest.c_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _07416_ (.A0(\sha256cu.m_out_digest.g_in[1] ),
    .A1(\sha256cu.m_out_digest.f_in[1] ),
    .S(\sha256cu.m_out_digest.e_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02045_));
 sky130_fd_sc_hd__and3_1 _07417_ (.A(_02043_),
    .B(_02044_),
    .C(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02046_));
 sky130_fd_sc_hd__a21o_1 _07418_ (.A1(_02043_),
    .A2(_02044_),
    .B1(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02047_));
 sky130_fd_sc_hd__and2b_1 _07419_ (.A_N(_02046_),
    .B(_02047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02048_));
 sky130_fd_sc_hd__xnor2_1 _07420_ (.A(\sha256cu.iter_processing.w[1] ),
    .B(_02048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02049_));
 sky130_fd_sc_hd__xnor2_1 _07421_ (.A(\sha256cu.m_out_digest.e_in[12] ),
    .B(\sha256cu.m_out_digest.e_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02050_));
 sky130_fd_sc_hd__xnor2_2 _07422_ (.A(\sha256cu.m_out_digest.e_in[26] ),
    .B(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02051_));
 sky130_fd_sc_hd__inv_2 _07423_ (.A(_02051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02052_));
 sky130_fd_sc_hd__xnor2_1 _07424_ (.A(\sha256cu.m_out_digest.a_in[14] ),
    .B(\sha256cu.m_out_digest.a_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02053_));
 sky130_fd_sc_hd__xnor2_2 _07425_ (.A(\sha256cu.m_out_digest.a_in[23] ),
    .B(_02053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02054_));
 sky130_fd_sc_hd__xnor2_1 _07426_ (.A(\sha256cu.m_out_digest.h_in[1] ),
    .B(_02054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02055_));
 sky130_fd_sc_hd__xnor2_1 _07427_ (.A(_02052_),
    .B(_02055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02056_));
 sky130_fd_sc_hd__nand2_1 _07428_ (.A(\sha256cu.m_out_digest.h_in[0] ),
    .B(_02029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02057_));
 sky130_fd_sc_hd__o21a_1 _07429_ (.A1(_02025_),
    .A2(_02030_),
    .B1(_02057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02058_));
 sky130_fd_sc_hd__xnor2_1 _07430_ (.A(_02056_),
    .B(_02058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02059_));
 sky130_fd_sc_hd__xor2_1 _07431_ (.A(_02049_),
    .B(_02059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02060_));
 sky130_fd_sc_hd__xnor2_1 _07432_ (.A(_02032_),
    .B(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02061_));
 sky130_fd_sc_hd__xnor2_1 _07433_ (.A(_02042_),
    .B(_02061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02062_));
 sky130_fd_sc_hd__xnor2_1 _07434_ (.A(\sha256cu.K[1] ),
    .B(_02062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_4 _07435_ (.A(_02005_),
    .B(_02015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_8 _07436_ (.A(_01911_),
    .B(_02064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02065_));
 sky130_fd_sc_hd__a21oi_1 _07437_ (.A1(_02035_),
    .A2(_02063_),
    .B1(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02066_));
 sky130_fd_sc_hd__o21a_1 _07438_ (.A1(_02035_),
    .A2(_02063_),
    .B1(_02066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02067_));
 sky130_fd_sc_hd__buf_6 _07439_ (.A(_02002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02068_));
 sky130_fd_sc_hd__a211o_1 _07440_ (.A1(\sha256cu.m_out_digest.a_in[1] ),
    .A2(_02040_),
    .B1(_02067_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00096_));
 sky130_fd_sc_hd__buf_6 _07441_ (.A(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02069_));
 sky130_fd_sc_hd__buf_4 _07442_ (.A(_02069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02070_));
 sky130_fd_sc_hd__inv_2 _07443_ (.A(\sha256cu.K[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02071_));
 sky130_fd_sc_hd__a21o_1 _07444_ (.A1(\sha256cu.iter_processing.w[1] ),
    .A2(_02047_),
    .B1(_02046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02072_));
 sky130_fd_sc_hd__or2_1 _07445_ (.A(\sha256cu.m_out_digest.b_in[2] ),
    .B(\sha256cu.m_out_digest.a_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02073_));
 sky130_fd_sc_hd__a21o_1 _07446_ (.A1(\sha256cu.m_out_digest.b_in[2] ),
    .A2(\sha256cu.m_out_digest.a_in[2] ),
    .B1(\sha256cu.m_out_digest.c_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _07447_ (.A0(\sha256cu.m_out_digest.g_in[2] ),
    .A1(\sha256cu.m_out_digest.f_in[2] ),
    .S(\sha256cu.m_out_digest.e_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02075_));
 sky130_fd_sc_hd__and3_1 _07448_ (.A(_02073_),
    .B(_02074_),
    .C(_02075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02076_));
 sky130_fd_sc_hd__a21o_1 _07449_ (.A1(_02073_),
    .A2(_02074_),
    .B1(_02075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02077_));
 sky130_fd_sc_hd__and2b_1 _07450_ (.A_N(_02076_),
    .B(_02077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02078_));
 sky130_fd_sc_hd__xnor2_1 _07451_ (.A(\sha256cu.iter_processing.w[2] ),
    .B(_02078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _07452_ (.A(\sha256cu.m_out_digest.e_in[13] ),
    .B(\sha256cu.m_out_digest.e_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02080_));
 sky130_fd_sc_hd__xnor2_2 _07453_ (.A(\sha256cu.m_out_digest.e_in[27] ),
    .B(_02080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02081_));
 sky130_fd_sc_hd__inv_2 _07454_ (.A(_02081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02082_));
 sky130_fd_sc_hd__buf_4 _07455_ (.A(\sha256cu.m_out_digest.a_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02083_));
 sky130_fd_sc_hd__clkbuf_4 _07456_ (.A(\sha256cu.m_out_digest.a_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02084_));
 sky130_fd_sc_hd__xnor2_1 _07457_ (.A(_02084_),
    .B(\sha256cu.m_out_digest.a_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02085_));
 sky130_fd_sc_hd__xnor2_1 _07458_ (.A(_02083_),
    .B(_02085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02086_));
 sky130_fd_sc_hd__xnor2_1 _07459_ (.A(\sha256cu.m_out_digest.h_in[2] ),
    .B(_02086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02087_));
 sky130_fd_sc_hd__xnor2_1 _07460_ (.A(_02082_),
    .B(_02087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2_1 _07461_ (.A(\sha256cu.m_out_digest.h_in[1] ),
    .B(_02054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02089_));
 sky130_fd_sc_hd__o21a_1 _07462_ (.A1(_02052_),
    .A2(_02055_),
    .B1(_02089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02090_));
 sky130_fd_sc_hd__xnor2_1 _07463_ (.A(_02088_),
    .B(_02090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02091_));
 sky130_fd_sc_hd__xor2_1 _07464_ (.A(_02079_),
    .B(_02091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_1 _07465_ (.A(_02056_),
    .B(_02058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02093_));
 sky130_fd_sc_hd__o21ba_1 _07466_ (.A1(_02049_),
    .A2(_02059_),
    .B1_N(_02093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02094_));
 sky130_fd_sc_hd__xnor2_1 _07467_ (.A(_02092_),
    .B(_02094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02095_));
 sky130_fd_sc_hd__xnor2_1 _07468_ (.A(_02072_),
    .B(_02095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02096_));
 sky130_fd_sc_hd__or2_1 _07469_ (.A(_02032_),
    .B(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02097_));
 sky130_fd_sc_hd__and2_1 _07470_ (.A(_02032_),
    .B(_02060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02098_));
 sky130_fd_sc_hd__a21oi_1 _07471_ (.A1(_02042_),
    .A2(_02097_),
    .B1(_02098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02099_));
 sky130_fd_sc_hd__xor2_1 _07472_ (.A(_02096_),
    .B(_02099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02100_));
 sky130_fd_sc_hd__xnor2_1 _07473_ (.A(_02071_),
    .B(_02100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02101_));
 sky130_fd_sc_hd__nand2_1 _07474_ (.A(\sha256cu.K[1] ),
    .B(_02062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02102_));
 sky130_fd_sc_hd__o21ai_1 _07475_ (.A1(_02035_),
    .A2(_02063_),
    .B1(_02102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02103_));
 sky130_fd_sc_hd__and2_1 _07476_ (.A(_02101_),
    .B(_02103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02104_));
 sky130_fd_sc_hd__nor2_1 _07477_ (.A(_02101_),
    .B(_02103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02105_));
 sky130_fd_sc_hd__or2_1 _07478_ (.A(_02104_),
    .B(_02105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02106_));
 sky130_fd_sc_hd__or2_1 _07479_ (.A(\sha256cu.m_out_digest.a_in[2] ),
    .B(_02002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02107_));
 sky130_fd_sc_hd__nand2_2 _07480_ (.A(_01564_),
    .B(_02064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02108_));
 sky130_fd_sc_hd__buf_2 _07481_ (.A(_02108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02109_));
 sky130_fd_sc_hd__buf_4 _07482_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02110_));
 sky130_fd_sc_hd__a2bb2o_1 _07483_ (.A1_N(_02070_),
    .A2_N(_02106_),
    .B1(_02107_),
    .B2(_02110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00097_));
 sky130_fd_sc_hd__clkbuf_8 _07484_ (.A(_01911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02111_));
 sky130_fd_sc_hd__nor2_4 _07485_ (.A(_02111_),
    .B(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02112_));
 sky130_fd_sc_hd__buf_4 _07486_ (.A(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02113_));
 sky130_fd_sc_hd__buf_4 _07487_ (.A(_02113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02114_));
 sky130_fd_sc_hd__or2_1 _07488_ (.A(_02096_),
    .B(_02099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02115_));
 sky130_fd_sc_hd__nand2_1 _07489_ (.A(\sha256cu.K[2] ),
    .B(_02100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02116_));
 sky130_fd_sc_hd__a21o_1 _07490_ (.A1(\sha256cu.iter_processing.w[2] ),
    .A2(_02077_),
    .B1(_02076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02117_));
 sky130_fd_sc_hd__or2_1 _07491_ (.A(\sha256cu.m_out_digest.b_in[3] ),
    .B(\sha256cu.m_out_digest.a_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02118_));
 sky130_fd_sc_hd__a21o_1 _07492_ (.A1(\sha256cu.m_out_digest.b_in[3] ),
    .A2(\sha256cu.m_out_digest.a_in[3] ),
    .B1(\sha256cu.m_out_digest.c_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _07493_ (.A0(\sha256cu.m_out_digest.g_in[3] ),
    .A1(\sha256cu.m_out_digest.f_in[3] ),
    .S(\sha256cu.m_out_digest.e_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02120_));
 sky130_fd_sc_hd__and3_1 _07494_ (.A(_02118_),
    .B(_02119_),
    .C(_02120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02121_));
 sky130_fd_sc_hd__a21o_1 _07495_ (.A1(_02118_),
    .A2(_02119_),
    .B1(_02120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02122_));
 sky130_fd_sc_hd__and2b_1 _07496_ (.A_N(_02121_),
    .B(_02122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02123_));
 sky130_fd_sc_hd__xnor2_1 _07497_ (.A(\sha256cu.iter_processing.w[3] ),
    .B(_02123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02124_));
 sky130_fd_sc_hd__xnor2_1 _07498_ (.A(\sha256cu.m_out_digest.e_in[14] ),
    .B(\sha256cu.m_out_digest.e_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02125_));
 sky130_fd_sc_hd__xnor2_2 _07499_ (.A(\sha256cu.m_out_digest.e_in[28] ),
    .B(_02125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02126_));
 sky130_fd_sc_hd__inv_2 _07500_ (.A(_02126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02127_));
 sky130_fd_sc_hd__clkbuf_4 _07501_ (.A(\sha256cu.m_out_digest.a_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02128_));
 sky130_fd_sc_hd__xnor2_1 _07502_ (.A(_02128_),
    .B(\sha256cu.m_out_digest.a_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02129_));
 sky130_fd_sc_hd__xnor2_1 _07503_ (.A(\sha256cu.m_out_digest.a_in[25] ),
    .B(_02129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02130_));
 sky130_fd_sc_hd__xnor2_1 _07504_ (.A(\sha256cu.m_out_digest.h_in[3] ),
    .B(_02130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02131_));
 sky130_fd_sc_hd__xnor2_1 _07505_ (.A(_02127_),
    .B(_02131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _07506_ (.A(\sha256cu.m_out_digest.h_in[2] ),
    .B(_02086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02133_));
 sky130_fd_sc_hd__o21a_1 _07507_ (.A1(_02082_),
    .A2(_02087_),
    .B1(_02133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02134_));
 sky130_fd_sc_hd__xnor2_1 _07508_ (.A(_02132_),
    .B(_02134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02135_));
 sky130_fd_sc_hd__xor2_1 _07509_ (.A(_02124_),
    .B(_02135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02136_));
 sky130_fd_sc_hd__nor2_1 _07510_ (.A(_02088_),
    .B(_02090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02137_));
 sky130_fd_sc_hd__o21ba_1 _07511_ (.A1(_02079_),
    .A2(_02091_),
    .B1_N(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02138_));
 sky130_fd_sc_hd__xnor2_1 _07512_ (.A(_02136_),
    .B(_02138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02139_));
 sky130_fd_sc_hd__xnor2_2 _07513_ (.A(_02117_),
    .B(_02139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02140_));
 sky130_fd_sc_hd__and2b_1 _07514_ (.A_N(_02094_),
    .B(_02092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02141_));
 sky130_fd_sc_hd__a21oi_2 _07515_ (.A1(_02072_),
    .A2(_02095_),
    .B1(_02141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02142_));
 sky130_fd_sc_hd__xor2_2 _07516_ (.A(_02140_),
    .B(_02142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02143_));
 sky130_fd_sc_hd__xnor2_1 _07517_ (.A(\sha256cu.K[3] ),
    .B(_02143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02144_));
 sky130_fd_sc_hd__nand3_1 _07518_ (.A(_02115_),
    .B(_02116_),
    .C(_02144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02145_));
 sky130_fd_sc_hd__a21oi_2 _07519_ (.A1(_02115_),
    .A2(_02116_),
    .B1(_02144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02146_));
 sky130_fd_sc_hd__inv_2 _07520_ (.A(_02146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_1 _07521_ (.A(_02145_),
    .B(_02147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02148_));
 sky130_fd_sc_hd__xnor2_1 _07522_ (.A(_02104_),
    .B(_02148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02149_));
 sky130_fd_sc_hd__a22o_1 _07523_ (.A1(\sha256cu.m_out_digest.a_in[3] ),
    .A2(_02070_),
    .B1(_02114_),
    .B2(_02149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00098_));
 sky130_fd_sc_hd__a21o_1 _07524_ (.A1(\sha256cu.iter_processing.w[3] ),
    .A2(_02122_),
    .B1(_02121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02150_));
 sky130_fd_sc_hd__or2_1 _07525_ (.A(\sha256cu.m_out_digest.b_in[4] ),
    .B(\sha256cu.m_out_digest.a_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02151_));
 sky130_fd_sc_hd__a21o_1 _07526_ (.A1(\sha256cu.m_out_digest.b_in[4] ),
    .A2(\sha256cu.m_out_digest.a_in[4] ),
    .B1(\sha256cu.m_out_digest.c_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02152_));
 sky130_fd_sc_hd__mux2_1 _07527_ (.A0(\sha256cu.m_out_digest.g_in[4] ),
    .A1(\sha256cu.m_out_digest.f_in[4] ),
    .S(\sha256cu.m_out_digest.e_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02153_));
 sky130_fd_sc_hd__and3_1 _07528_ (.A(_02151_),
    .B(_02152_),
    .C(_02153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02154_));
 sky130_fd_sc_hd__a21o_1 _07529_ (.A1(_02151_),
    .A2(_02152_),
    .B1(_02153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02155_));
 sky130_fd_sc_hd__and2b_1 _07530_ (.A_N(_02154_),
    .B(_02155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02156_));
 sky130_fd_sc_hd__xnor2_1 _07531_ (.A(\sha256cu.iter_processing.w[4] ),
    .B(_02156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_1 _07532_ (.A(\sha256cu.m_out_digest.e_in[15] ),
    .B(\sha256cu.m_out_digest.e_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02158_));
 sky130_fd_sc_hd__xnor2_2 _07533_ (.A(\sha256cu.m_out_digest.e_in[29] ),
    .B(_02158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02159_));
 sky130_fd_sc_hd__inv_2 _07534_ (.A(_02159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02160_));
 sky130_fd_sc_hd__buf_4 _07535_ (.A(\sha256cu.m_out_digest.a_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02161_));
 sky130_fd_sc_hd__clkbuf_4 _07536_ (.A(\sha256cu.m_out_digest.a_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02162_));
 sky130_fd_sc_hd__xnor2_1 _07537_ (.A(_02162_),
    .B(\sha256cu.m_out_digest.a_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02163_));
 sky130_fd_sc_hd__xnor2_1 _07538_ (.A(_02161_),
    .B(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02164_));
 sky130_fd_sc_hd__xnor2_1 _07539_ (.A(\sha256cu.m_out_digest.h_in[4] ),
    .B(_02164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_1 _07540_ (.A(_02160_),
    .B(_02165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02166_));
 sky130_fd_sc_hd__nand2_1 _07541_ (.A(\sha256cu.m_out_digest.h_in[3] ),
    .B(_02130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02167_));
 sky130_fd_sc_hd__o21a_1 _07542_ (.A1(_02127_),
    .A2(_02131_),
    .B1(_02167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02168_));
 sky130_fd_sc_hd__xnor2_1 _07543_ (.A(_02166_),
    .B(_02168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02169_));
 sky130_fd_sc_hd__xor2_1 _07544_ (.A(_02157_),
    .B(_02169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02170_));
 sky130_fd_sc_hd__nor2_1 _07545_ (.A(_02132_),
    .B(_02134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02171_));
 sky130_fd_sc_hd__o21ba_1 _07546_ (.A1(_02124_),
    .A2(_02135_),
    .B1_N(_02171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02172_));
 sky130_fd_sc_hd__xnor2_1 _07547_ (.A(_02170_),
    .B(_02172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02173_));
 sky130_fd_sc_hd__xnor2_1 _07548_ (.A(_02150_),
    .B(_02173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02174_));
 sky130_fd_sc_hd__and2b_1 _07549_ (.A_N(_02138_),
    .B(_02136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02175_));
 sky130_fd_sc_hd__a21oi_1 _07550_ (.A1(_02117_),
    .A2(_02139_),
    .B1(_02175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02176_));
 sky130_fd_sc_hd__xor2_1 _07551_ (.A(_02174_),
    .B(_02176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02177_));
 sky130_fd_sc_hd__xnor2_1 _07552_ (.A(\sha256cu.K[4] ),
    .B(_02177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _07553_ (.A(_02140_),
    .B(_02142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02179_));
 sky130_fd_sc_hd__a21oi_2 _07554_ (.A1(\sha256cu.K[3] ),
    .A2(_02143_),
    .B1(_02179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02180_));
 sky130_fd_sc_hd__xor2_1 _07555_ (.A(_02178_),
    .B(_02180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02181_));
 sky130_fd_sc_hd__o21a_1 _07556_ (.A1(_02104_),
    .A2(_02146_),
    .B1(_02145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02182_));
 sky130_fd_sc_hd__nand2_1 _07557_ (.A(_02181_),
    .B(_02182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02183_));
 sky130_fd_sc_hd__o21a_1 _07558_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02184_));
 sky130_fd_sc_hd__a22o_1 _07559_ (.A1(\sha256cu.m_out_digest.a_in[4] ),
    .A2(_02070_),
    .B1(_02183_),
    .B2(_02184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00099_));
 sky130_fd_sc_hd__nor2_1 _07560_ (.A(_02174_),
    .B(_02176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02185_));
 sky130_fd_sc_hd__a21oi_1 _07561_ (.A1(\sha256cu.K[4] ),
    .A2(_02177_),
    .B1(_02185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02186_));
 sky130_fd_sc_hd__a21o_1 _07562_ (.A1(\sha256cu.iter_processing.w[4] ),
    .A2(_02155_),
    .B1(_02154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02187_));
 sky130_fd_sc_hd__or2_1 _07563_ (.A(\sha256cu.m_out_digest.b_in[5] ),
    .B(\sha256cu.m_out_digest.a_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02188_));
 sky130_fd_sc_hd__a21o_1 _07564_ (.A1(\sha256cu.m_out_digest.b_in[5] ),
    .A2(\sha256cu.m_out_digest.a_in[5] ),
    .B1(\sha256cu.m_out_digest.c_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _07565_ (.A0(\sha256cu.m_out_digest.g_in[5] ),
    .A1(\sha256cu.m_out_digest.f_in[5] ),
    .S(\sha256cu.m_out_digest.e_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02190_));
 sky130_fd_sc_hd__and3_1 _07566_ (.A(_02188_),
    .B(_02189_),
    .C(_02190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02191_));
 sky130_fd_sc_hd__a21o_1 _07567_ (.A1(_02188_),
    .A2(_02189_),
    .B1(_02190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02192_));
 sky130_fd_sc_hd__and2b_1 _07568_ (.A_N(_02191_),
    .B(_02192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_1 _07569_ (.A(\sha256cu.iter_processing.w[5] ),
    .B(_02193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02194_));
 sky130_fd_sc_hd__xnor2_2 _07570_ (.A(\sha256cu.m_out_digest.e_in[16] ),
    .B(\sha256cu.m_out_digest.e_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02195_));
 sky130_fd_sc_hd__xnor2_4 _07571_ (.A(\sha256cu.m_out_digest.e_in[30] ),
    .B(_02195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02196_));
 sky130_fd_sc_hd__inv_2 _07572_ (.A(_02196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02197_));
 sky130_fd_sc_hd__clkbuf_4 _07573_ (.A(\sha256cu.m_out_digest.a_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02198_));
 sky130_fd_sc_hd__xnor2_1 _07574_ (.A(_02198_),
    .B(\sha256cu.m_out_digest.a_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _07575_ (.A(\sha256cu.m_out_digest.a_in[27] ),
    .B(_02199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02200_));
 sky130_fd_sc_hd__xnor2_1 _07576_ (.A(\sha256cu.m_out_digest.h_in[5] ),
    .B(_02200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02201_));
 sky130_fd_sc_hd__xnor2_1 _07577_ (.A(_02197_),
    .B(_02201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02202_));
 sky130_fd_sc_hd__nand2_1 _07578_ (.A(\sha256cu.m_out_digest.h_in[4] ),
    .B(_02164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02203_));
 sky130_fd_sc_hd__o21a_1 _07579_ (.A1(_02160_),
    .A2(_02165_),
    .B1(_02203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02204_));
 sky130_fd_sc_hd__xnor2_1 _07580_ (.A(_02202_),
    .B(_02204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02205_));
 sky130_fd_sc_hd__xor2_1 _07581_ (.A(_02194_),
    .B(_02205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02206_));
 sky130_fd_sc_hd__nor2_1 _07582_ (.A(_02166_),
    .B(_02168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02207_));
 sky130_fd_sc_hd__o21ba_1 _07583_ (.A1(_02157_),
    .A2(_02169_),
    .B1_N(_02207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02208_));
 sky130_fd_sc_hd__xnor2_1 _07584_ (.A(_02206_),
    .B(_02208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02209_));
 sky130_fd_sc_hd__xnor2_1 _07585_ (.A(_02187_),
    .B(_02209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02210_));
 sky130_fd_sc_hd__and2b_1 _07586_ (.A_N(_02172_),
    .B(_02170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02211_));
 sky130_fd_sc_hd__a21oi_1 _07587_ (.A1(_02150_),
    .A2(_02173_),
    .B1(_02211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02212_));
 sky130_fd_sc_hd__xor2_1 _07588_ (.A(_02210_),
    .B(_02212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02213_));
 sky130_fd_sc_hd__xnor2_1 _07589_ (.A(\sha256cu.K[5] ),
    .B(_02213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02214_));
 sky130_fd_sc_hd__xor2_1 _07590_ (.A(_02186_),
    .B(_02214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02215_));
 sky130_fd_sc_hd__o21a_1 _07591_ (.A1(_02178_),
    .A2(_02180_),
    .B1(_02183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02216_));
 sky130_fd_sc_hd__xnor2_1 _07592_ (.A(_02215_),
    .B(_02216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02217_));
 sky130_fd_sc_hd__a22o_1 _07593_ (.A1(\sha256cu.m_out_digest.a_in[5] ),
    .A2(_02037_),
    .B1(_02017_),
    .B2(_02217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02218_));
 sky130_fd_sc_hd__or2_1 _07594_ (.A(_01913_),
    .B(_02218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02219_));
 sky130_fd_sc_hd__clkbuf_1 _07595_ (.A(_02219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00100_));
 sky130_fd_sc_hd__clkbuf_8 _07596_ (.A(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02220_));
 sky130_fd_sc_hd__a21o_1 _07597_ (.A1(\sha256cu.iter_processing.w[5] ),
    .A2(_02192_),
    .B1(_02191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02221_));
 sky130_fd_sc_hd__or2_1 _07598_ (.A(\sha256cu.m_out_digest.b_in[6] ),
    .B(\sha256cu.m_out_digest.a_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02222_));
 sky130_fd_sc_hd__a21o_1 _07599_ (.A1(\sha256cu.m_out_digest.b_in[6] ),
    .A2(\sha256cu.m_out_digest.a_in[6] ),
    .B1(\sha256cu.m_out_digest.c_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _07600_ (.A0(\sha256cu.m_out_digest.g_in[6] ),
    .A1(\sha256cu.m_out_digest.f_in[6] ),
    .S(\sha256cu.m_out_digest.e_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02224_));
 sky130_fd_sc_hd__and3_1 _07601_ (.A(_02222_),
    .B(_02223_),
    .C(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02225_));
 sky130_fd_sc_hd__a21o_1 _07602_ (.A1(_02222_),
    .A2(_02223_),
    .B1(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02226_));
 sky130_fd_sc_hd__and2b_1 _07603_ (.A_N(_02225_),
    .B(_02226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02227_));
 sky130_fd_sc_hd__xnor2_2 _07604_ (.A(\sha256cu.iter_processing.w[6] ),
    .B(_02227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02228_));
 sky130_fd_sc_hd__xnor2_1 _07605_ (.A(\sha256cu.m_out_digest.e_in[17] ),
    .B(\sha256cu.m_out_digest.e_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02229_));
 sky130_fd_sc_hd__xnor2_2 _07606_ (.A(\sha256cu.m_out_digest.e_in[31] ),
    .B(_02229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02230_));
 sky130_fd_sc_hd__inv_2 _07607_ (.A(_02230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02231_));
 sky130_fd_sc_hd__buf_4 _07608_ (.A(\sha256cu.m_out_digest.a_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_4 _07609_ (.A(\sha256cu.m_out_digest.a_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02233_));
 sky130_fd_sc_hd__xnor2_2 _07610_ (.A(_02233_),
    .B(\sha256cu.m_out_digest.a_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02234_));
 sky130_fd_sc_hd__xnor2_4 _07611_ (.A(_02232_),
    .B(_02234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02235_));
 sky130_fd_sc_hd__xnor2_2 _07612_ (.A(\sha256cu.m_out_digest.h_in[6] ),
    .B(_02235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02236_));
 sky130_fd_sc_hd__xnor2_2 _07613_ (.A(_02231_),
    .B(_02236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_1 _07614_ (.A(\sha256cu.m_out_digest.h_in[5] ),
    .B(_02200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02238_));
 sky130_fd_sc_hd__o21a_1 _07615_ (.A1(_02197_),
    .A2(_02201_),
    .B1(_02238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02239_));
 sky130_fd_sc_hd__xnor2_2 _07616_ (.A(_02237_),
    .B(_02239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02240_));
 sky130_fd_sc_hd__xor2_2 _07617_ (.A(_02228_),
    .B(_02240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02241_));
 sky130_fd_sc_hd__nor2_1 _07618_ (.A(_02202_),
    .B(_02204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02242_));
 sky130_fd_sc_hd__o21ba_1 _07619_ (.A1(_02194_),
    .A2(_02205_),
    .B1_N(_02242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02243_));
 sky130_fd_sc_hd__xnor2_2 _07620_ (.A(_02241_),
    .B(_02243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02244_));
 sky130_fd_sc_hd__xnor2_2 _07621_ (.A(_02221_),
    .B(_02244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02245_));
 sky130_fd_sc_hd__or2b_1 _07622_ (.A(_02208_),
    .B_N(_02206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02246_));
 sky130_fd_sc_hd__a21boi_2 _07623_ (.A1(_02187_),
    .A2(_02209_),
    .B1_N(_02246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02247_));
 sky130_fd_sc_hd__xor2_2 _07624_ (.A(_02245_),
    .B(_02247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02248_));
 sky130_fd_sc_hd__xnor2_2 _07625_ (.A(\sha256cu.K[6] ),
    .B(_02248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02249_));
 sky130_fd_sc_hd__nor2_1 _07626_ (.A(_02210_),
    .B(_02212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02250_));
 sky130_fd_sc_hd__a21oi_2 _07627_ (.A1(\sha256cu.K[5] ),
    .A2(_02213_),
    .B1(_02250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02251_));
 sky130_fd_sc_hd__xnor2_2 _07628_ (.A(_02249_),
    .B(_02251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02252_));
 sky130_fd_sc_hd__o22a_1 _07629_ (.A1(_02178_),
    .A2(_02180_),
    .B1(_02186_),
    .B2(_02214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02253_));
 sky130_fd_sc_hd__and2_1 _07630_ (.A(_02186_),
    .B(_02214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02254_));
 sky130_fd_sc_hd__a21o_1 _07631_ (.A1(_02183_),
    .A2(_02253_),
    .B1(_02254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02255_));
 sky130_fd_sc_hd__or2_1 _07632_ (.A(_02252_),
    .B(_02255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02256_));
 sky130_fd_sc_hd__a21oi_1 _07633_ (.A1(_02252_),
    .A2(_02255_),
    .B1(_02069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02257_));
 sky130_fd_sc_hd__buf_4 _07634_ (.A(_02002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02258_));
 sky130_fd_sc_hd__a221o_1 _07635_ (.A1(\sha256cu.m_out_digest.a_in[6] ),
    .A2(_02220_),
    .B1(_02256_),
    .B2(_02257_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00101_));
 sky130_fd_sc_hd__nor2_1 _07636_ (.A(_02245_),
    .B(_02247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02259_));
 sky130_fd_sc_hd__a21oi_2 _07637_ (.A1(\sha256cu.K[6] ),
    .A2(_02248_),
    .B1(_02259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02260_));
 sky130_fd_sc_hd__a21o_1 _07638_ (.A1(\sha256cu.iter_processing.w[6] ),
    .A2(_02226_),
    .B1(_02225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02261_));
 sky130_fd_sc_hd__or2_1 _07639_ (.A(\sha256cu.m_out_digest.b_in[7] ),
    .B(\sha256cu.m_out_digest.a_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02262_));
 sky130_fd_sc_hd__a21o_1 _07640_ (.A1(\sha256cu.m_out_digest.b_in[7] ),
    .A2(\sha256cu.m_out_digest.a_in[7] ),
    .B1(\sha256cu.m_out_digest.c_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _07641_ (.A0(\sha256cu.m_out_digest.g_in[7] ),
    .A1(\sha256cu.m_out_digest.f_in[7] ),
    .S(\sha256cu.m_out_digest.e_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02264_));
 sky130_fd_sc_hd__and3_1 _07642_ (.A(_02262_),
    .B(_02263_),
    .C(_02264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02265_));
 sky130_fd_sc_hd__a21o_1 _07643_ (.A1(_02262_),
    .A2(_02263_),
    .B1(_02264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02266_));
 sky130_fd_sc_hd__and2b_1 _07644_ (.A_N(_02265_),
    .B(_02266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02267_));
 sky130_fd_sc_hd__xnor2_2 _07645_ (.A(\sha256cu.iter_processing.w[7] ),
    .B(_02267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02268_));
 sky130_fd_sc_hd__xnor2_1 _07646_ (.A(\sha256cu.m_out_digest.e_in[13] ),
    .B(\sha256cu.m_out_digest.e_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02269_));
 sky130_fd_sc_hd__xnor2_2 _07647_ (.A(\sha256cu.m_out_digest.e_in[18] ),
    .B(_02269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02270_));
 sky130_fd_sc_hd__inv_2 _07648_ (.A(_02270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02271_));
 sky130_fd_sc_hd__buf_4 _07649_ (.A(\sha256cu.m_out_digest.a_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02272_));
 sky130_fd_sc_hd__buf_4 _07650_ (.A(\sha256cu.m_out_digest.a_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02273_));
 sky130_fd_sc_hd__xnor2_4 _07651_ (.A(_02273_),
    .B(\sha256cu.m_out_digest.a_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02274_));
 sky130_fd_sc_hd__xnor2_4 _07652_ (.A(_02272_),
    .B(_02274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02275_));
 sky130_fd_sc_hd__xnor2_2 _07653_ (.A(\sha256cu.m_out_digest.h_in[7] ),
    .B(_02275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02276_));
 sky130_fd_sc_hd__xnor2_2 _07654_ (.A(_02271_),
    .B(_02276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _07655_ (.A(\sha256cu.m_out_digest.h_in[6] ),
    .B(_02235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02278_));
 sky130_fd_sc_hd__o21a_1 _07656_ (.A1(_02231_),
    .A2(_02236_),
    .B1(_02278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02279_));
 sky130_fd_sc_hd__xnor2_2 _07657_ (.A(_02277_),
    .B(_02279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02280_));
 sky130_fd_sc_hd__xor2_2 _07658_ (.A(_02268_),
    .B(_02280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02281_));
 sky130_fd_sc_hd__nor2_1 _07659_ (.A(_02237_),
    .B(_02239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02282_));
 sky130_fd_sc_hd__o21ba_1 _07660_ (.A1(_02228_),
    .A2(_02240_),
    .B1_N(_02282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02283_));
 sky130_fd_sc_hd__xnor2_2 _07661_ (.A(_02281_),
    .B(_02283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02284_));
 sky130_fd_sc_hd__xnor2_2 _07662_ (.A(_02261_),
    .B(_02284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02285_));
 sky130_fd_sc_hd__and2b_1 _07663_ (.A_N(_02243_),
    .B(_02241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02286_));
 sky130_fd_sc_hd__a21oi_2 _07664_ (.A1(_02221_),
    .A2(_02244_),
    .B1(_02286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02287_));
 sky130_fd_sc_hd__xor2_2 _07665_ (.A(_02285_),
    .B(_02287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02288_));
 sky130_fd_sc_hd__xnor2_2 _07666_ (.A(\sha256cu.K[7] ),
    .B(_02288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02289_));
 sky130_fd_sc_hd__xnor2_2 _07667_ (.A(_02260_),
    .B(_02289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02290_));
 sky130_fd_sc_hd__o21ai_1 _07668_ (.A1(_02249_),
    .A2(_02251_),
    .B1(_02256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02291_));
 sky130_fd_sc_hd__xnor2_1 _07669_ (.A(_02290_),
    .B(_02291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02292_));
 sky130_fd_sc_hd__a22o_1 _07670_ (.A1(\sha256cu.m_out_digest.a_in[7] ),
    .A2(_02070_),
    .B1(_02114_),
    .B2(_02292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00102_));
 sky130_fd_sc_hd__a21o_1 _07671_ (.A1(\sha256cu.iter_processing.w[7] ),
    .A2(_02266_),
    .B1(_02265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02293_));
 sky130_fd_sc_hd__or2_1 _07672_ (.A(\sha256cu.m_out_digest.b_in[8] ),
    .B(\sha256cu.m_out_digest.a_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02294_));
 sky130_fd_sc_hd__a21o_1 _07673_ (.A1(\sha256cu.m_out_digest.b_in[8] ),
    .A2(\sha256cu.m_out_digest.a_in[8] ),
    .B1(\sha256cu.m_out_digest.c_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _07674_ (.A0(\sha256cu.m_out_digest.g_in[8] ),
    .A1(\sha256cu.m_out_digest.f_in[8] ),
    .S(\sha256cu.m_out_digest.e_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02296_));
 sky130_fd_sc_hd__and3_1 _07675_ (.A(_02294_),
    .B(_02295_),
    .C(_02296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02297_));
 sky130_fd_sc_hd__a21o_1 _07676_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02298_));
 sky130_fd_sc_hd__and2b_1 _07677_ (.A_N(_02297_),
    .B(_02298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02299_));
 sky130_fd_sc_hd__xnor2_2 _07678_ (.A(\sha256cu.iter_processing.w[8] ),
    .B(_02299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02300_));
 sky130_fd_sc_hd__xnor2_2 _07679_ (.A(\sha256cu.m_out_digest.e_in[14] ),
    .B(\sha256cu.m_out_digest.e_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02301_));
 sky130_fd_sc_hd__xnor2_4 _07680_ (.A(\sha256cu.m_out_digest.e_in[19] ),
    .B(_02301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02302_));
 sky130_fd_sc_hd__inv_2 _07681_ (.A(_02302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02303_));
 sky130_fd_sc_hd__buf_4 _07682_ (.A(\sha256cu.m_out_digest.a_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02304_));
 sky130_fd_sc_hd__xnor2_2 _07683_ (.A(\sha256cu.m_out_digest.a_in[21] ),
    .B(\sha256cu.m_out_digest.a_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02305_));
 sky130_fd_sc_hd__xnor2_4 _07684_ (.A(_02304_),
    .B(_02305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02306_));
 sky130_fd_sc_hd__xnor2_2 _07685_ (.A(\sha256cu.m_out_digest.h_in[8] ),
    .B(_02306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02307_));
 sky130_fd_sc_hd__xnor2_2 _07686_ (.A(_02303_),
    .B(_02307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02308_));
 sky130_fd_sc_hd__nand2_1 _07687_ (.A(\sha256cu.m_out_digest.h_in[7] ),
    .B(_02275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02309_));
 sky130_fd_sc_hd__o21a_1 _07688_ (.A1(_02271_),
    .A2(_02276_),
    .B1(_02309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02310_));
 sky130_fd_sc_hd__xnor2_2 _07689_ (.A(_02308_),
    .B(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02311_));
 sky130_fd_sc_hd__xor2_2 _07690_ (.A(_02300_),
    .B(_02311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02312_));
 sky130_fd_sc_hd__nor2_1 _07691_ (.A(_02277_),
    .B(_02279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02313_));
 sky130_fd_sc_hd__o21ba_1 _07692_ (.A1(_02268_),
    .A2(_02280_),
    .B1_N(_02313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02314_));
 sky130_fd_sc_hd__xnor2_2 _07693_ (.A(_02312_),
    .B(_02314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02315_));
 sky130_fd_sc_hd__xnor2_2 _07694_ (.A(_02293_),
    .B(_02315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02316_));
 sky130_fd_sc_hd__or2b_1 _07695_ (.A(_02283_),
    .B_N(_02281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02317_));
 sky130_fd_sc_hd__a21bo_1 _07696_ (.A1(_02261_),
    .A2(_02284_),
    .B1_N(_02317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02318_));
 sky130_fd_sc_hd__xnor2_2 _07697_ (.A(_02316_),
    .B(_02318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02319_));
 sky130_fd_sc_hd__xnor2_2 _07698_ (.A(\sha256cu.K[8] ),
    .B(_02319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _07699_ (.A(_02285_),
    .B(_02287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02321_));
 sky130_fd_sc_hd__a21o_1 _07700_ (.A1(\sha256cu.K[7] ),
    .A2(_02288_),
    .B1(_02321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02322_));
 sky130_fd_sc_hd__xor2_2 _07701_ (.A(_02320_),
    .B(_02322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02323_));
 sky130_fd_sc_hd__o2111a_1 _07702_ (.A1(_02104_),
    .A2(_02146_),
    .B1(_02181_),
    .C1(_02215_),
    .D1(_02145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02324_));
 sky130_fd_sc_hd__nor2_1 _07703_ (.A(_02252_),
    .B(_02290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02325_));
 sky130_fd_sc_hd__nor4_2 _07704_ (.A(_02254_),
    .B(_02252_),
    .C(_02253_),
    .D(_02290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02326_));
 sky130_fd_sc_hd__a211o_1 _07705_ (.A1(_02260_),
    .A2(_02289_),
    .B1(_02249_),
    .C1(_02251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02327_));
 sky130_fd_sc_hd__o21ai_1 _07706_ (.A1(_02260_),
    .A2(_02289_),
    .B1(_02327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02328_));
 sky130_fd_sc_hd__a211oi_4 _07707_ (.A1(_02324_),
    .A2(_02325_),
    .B1(_02326_),
    .C1(_02328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _07708_ (.A(_02323_),
    .B(_02329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02330_));
 sky130_fd_sc_hd__or2_1 _07709_ (.A(_02323_),
    .B(_02329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02331_));
 sky130_fd_sc_hd__buf_4 _07710_ (.A(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02332_));
 sky130_fd_sc_hd__a32o_1 _07711_ (.A1(_02113_),
    .A2(_02330_),
    .A3(_02331_),
    .B1(_02332_),
    .B2(\sha256cu.m_out_digest.a_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00103_));
 sky130_fd_sc_hd__or2b_1 _07712_ (.A(_02316_),
    .B_N(_02318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02333_));
 sky130_fd_sc_hd__a21boi_1 _07713_ (.A1(\sha256cu.K[8] ),
    .A2(_02319_),
    .B1_N(_02333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02334_));
 sky130_fd_sc_hd__a21o_1 _07714_ (.A1(\sha256cu.iter_processing.w[8] ),
    .A2(_02298_),
    .B1(_02297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02335_));
 sky130_fd_sc_hd__or2_1 _07715_ (.A(\sha256cu.m_out_digest.b_in[9] ),
    .B(\sha256cu.m_out_digest.a_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02336_));
 sky130_fd_sc_hd__a21o_1 _07716_ (.A1(\sha256cu.m_out_digest.b_in[9] ),
    .A2(\sha256cu.m_out_digest.a_in[9] ),
    .B1(\sha256cu.m_out_digest.c_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02337_));
 sky130_fd_sc_hd__mux2_1 _07717_ (.A0(\sha256cu.m_out_digest.g_in[9] ),
    .A1(\sha256cu.m_out_digest.f_in[9] ),
    .S(\sha256cu.m_out_digest.e_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02338_));
 sky130_fd_sc_hd__and3_1 _07718_ (.A(_02336_),
    .B(_02337_),
    .C(_02338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02339_));
 sky130_fd_sc_hd__a21o_1 _07719_ (.A1(_02336_),
    .A2(_02337_),
    .B1(_02338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02340_));
 sky130_fd_sc_hd__and2b_1 _07720_ (.A_N(_02339_),
    .B(_02340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02341_));
 sky130_fd_sc_hd__xnor2_1 _07721_ (.A(\sha256cu.iter_processing.w[9] ),
    .B(_02341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02342_));
 sky130_fd_sc_hd__xnor2_2 _07722_ (.A(\sha256cu.m_out_digest.e_in[15] ),
    .B(\sha256cu.m_out_digest.e_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02343_));
 sky130_fd_sc_hd__xnor2_4 _07723_ (.A(\sha256cu.m_out_digest.e_in[20] ),
    .B(_02343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02344_));
 sky130_fd_sc_hd__inv_2 _07724_ (.A(_02344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02345_));
 sky130_fd_sc_hd__xnor2_2 _07725_ (.A(_02026_),
    .B(\sha256cu.m_out_digest.a_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02346_));
 sky130_fd_sc_hd__xnor2_4 _07726_ (.A(\sha256cu.m_out_digest.a_in[31] ),
    .B(_02346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02347_));
 sky130_fd_sc_hd__xnor2_1 _07727_ (.A(\sha256cu.m_out_digest.h_in[9] ),
    .B(_02347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02348_));
 sky130_fd_sc_hd__xnor2_1 _07728_ (.A(_02345_),
    .B(_02348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02349_));
 sky130_fd_sc_hd__nand2_1 _07729_ (.A(\sha256cu.m_out_digest.h_in[8] ),
    .B(_02306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02350_));
 sky130_fd_sc_hd__o21a_1 _07730_ (.A1(_02303_),
    .A2(_02307_),
    .B1(_02350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02351_));
 sky130_fd_sc_hd__xnor2_1 _07731_ (.A(_02349_),
    .B(_02351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02352_));
 sky130_fd_sc_hd__xor2_1 _07732_ (.A(_02342_),
    .B(_02352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02353_));
 sky130_fd_sc_hd__nor2_1 _07733_ (.A(_02308_),
    .B(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02354_));
 sky130_fd_sc_hd__o21ba_1 _07734_ (.A1(_02300_),
    .A2(_02311_),
    .B1_N(_02354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02355_));
 sky130_fd_sc_hd__xnor2_1 _07735_ (.A(_02353_),
    .B(_02355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02356_));
 sky130_fd_sc_hd__xnor2_1 _07736_ (.A(_02335_),
    .B(_02356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02357_));
 sky130_fd_sc_hd__and2b_1 _07737_ (.A_N(_02314_),
    .B(_02312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02358_));
 sky130_fd_sc_hd__a21oi_1 _07738_ (.A1(_02293_),
    .A2(_02315_),
    .B1(_02358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02359_));
 sky130_fd_sc_hd__xor2_1 _07739_ (.A(_02357_),
    .B(_02359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02360_));
 sky130_fd_sc_hd__xnor2_1 _07740_ (.A(\sha256cu.K[9] ),
    .B(_02360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_1 _07741_ (.A(_02334_),
    .B(_02361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02362_));
 sky130_fd_sc_hd__or2_1 _07742_ (.A(_02334_),
    .B(_02361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02363_));
 sky130_fd_sc_hd__nand2_1 _07743_ (.A(_02362_),
    .B(_02363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02364_));
 sky130_fd_sc_hd__and2b_1 _07744_ (.A_N(_02320_),
    .B(_02322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02365_));
 sky130_fd_sc_hd__o21ba_1 _07745_ (.A1(_02323_),
    .A2(_02329_),
    .B1_N(_02365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02366_));
 sky130_fd_sc_hd__xnor2_1 _07746_ (.A(_02364_),
    .B(_02366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_1 _07747_ (.A(_02069_),
    .B(_02367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02368_));
 sky130_fd_sc_hd__a211o_1 _07748_ (.A1(\sha256cu.m_out_digest.a_in[9] ),
    .A2(_02040_),
    .B1(_02368_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00104_));
 sky130_fd_sc_hd__clkbuf_4 _07749_ (.A(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02369_));
 sky130_fd_sc_hd__buf_4 _07750_ (.A(_02369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02370_));
 sky130_fd_sc_hd__a21o_1 _07751_ (.A1(\sha256cu.iter_processing.w[9] ),
    .A2(_02340_),
    .B1(_02339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02371_));
 sky130_fd_sc_hd__or2_1 _07752_ (.A(\sha256cu.m_out_digest.b_in[10] ),
    .B(\sha256cu.m_out_digest.a_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02372_));
 sky130_fd_sc_hd__a21o_1 _07753_ (.A1(\sha256cu.m_out_digest.b_in[10] ),
    .A2(\sha256cu.m_out_digest.a_in[10] ),
    .B1(\sha256cu.m_out_digest.c_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02373_));
 sky130_fd_sc_hd__mux2_1 _07754_ (.A0(\sha256cu.m_out_digest.g_in[10] ),
    .A1(\sha256cu.m_out_digest.f_in[10] ),
    .S(\sha256cu.m_out_digest.e_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02374_));
 sky130_fd_sc_hd__and3_1 _07755_ (.A(_02372_),
    .B(_02373_),
    .C(_02374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02375_));
 sky130_fd_sc_hd__a21o_1 _07756_ (.A1(_02372_),
    .A2(_02373_),
    .B1(_02374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02376_));
 sky130_fd_sc_hd__and2b_1 _07757_ (.A_N(_02375_),
    .B(_02376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02377_));
 sky130_fd_sc_hd__xnor2_1 _07758_ (.A(\sha256cu.iter_processing.w[10] ),
    .B(_02377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02378_));
 sky130_fd_sc_hd__xnor2_1 _07759_ (.A(\sha256cu.m_out_digest.e_in[16] ),
    .B(\sha256cu.m_out_digest.e_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02379_));
 sky130_fd_sc_hd__xnor2_2 _07760_ (.A(\sha256cu.m_out_digest.e_in[21] ),
    .B(_02379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02380_));
 sky130_fd_sc_hd__inv_2 _07761_ (.A(_02380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02381_));
 sky130_fd_sc_hd__clkbuf_4 _07762_ (.A(\sha256cu.m_out_digest.a_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02382_));
 sky130_fd_sc_hd__xnor2_1 _07763_ (.A(_02382_),
    .B(\sha256cu.m_out_digest.a_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02383_));
 sky130_fd_sc_hd__xnor2_2 _07764_ (.A(\sha256cu.m_out_digest.a_in[23] ),
    .B(_02383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02384_));
 sky130_fd_sc_hd__xnor2_1 _07765_ (.A(\sha256cu.m_out_digest.h_in[10] ),
    .B(_02384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02385_));
 sky130_fd_sc_hd__xnor2_1 _07766_ (.A(_02381_),
    .B(_02385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _07767_ (.A(\sha256cu.m_out_digest.h_in[9] ),
    .B(_02347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02387_));
 sky130_fd_sc_hd__o21a_1 _07768_ (.A1(_02345_),
    .A2(_02348_),
    .B1(_02387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02388_));
 sky130_fd_sc_hd__xnor2_1 _07769_ (.A(_02386_),
    .B(_02388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02389_));
 sky130_fd_sc_hd__xor2_1 _07770_ (.A(_02378_),
    .B(_02389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02390_));
 sky130_fd_sc_hd__nor2_1 _07771_ (.A(_02349_),
    .B(_02351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02391_));
 sky130_fd_sc_hd__o21ba_1 _07772_ (.A1(_02342_),
    .A2(_02352_),
    .B1_N(_02391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02392_));
 sky130_fd_sc_hd__xnor2_1 _07773_ (.A(_02390_),
    .B(_02392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02393_));
 sky130_fd_sc_hd__xnor2_1 _07774_ (.A(_02371_),
    .B(_02393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02394_));
 sky130_fd_sc_hd__or2b_1 _07775_ (.A(_02355_),
    .B_N(_02353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02395_));
 sky130_fd_sc_hd__a21bo_1 _07776_ (.A1(_02335_),
    .A2(_02356_),
    .B1_N(_02395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02396_));
 sky130_fd_sc_hd__xnor2_1 _07777_ (.A(_02394_),
    .B(_02396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02397_));
 sky130_fd_sc_hd__xnor2_1 _07778_ (.A(\sha256cu.K[10] ),
    .B(_02397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _07779_ (.A(_02357_),
    .B(_02359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02399_));
 sky130_fd_sc_hd__a21oi_1 _07780_ (.A1(\sha256cu.K[9] ),
    .A2(_02360_),
    .B1(_02399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02400_));
 sky130_fd_sc_hd__xnor2_1 _07781_ (.A(_02398_),
    .B(_02400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02401_));
 sky130_fd_sc_hd__and3b_1 _07782_ (.A_N(_02323_),
    .B(_02362_),
    .C(_02363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02402_));
 sky130_fd_sc_hd__inv_2 _07783_ (.A(_02402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _07784_ (.A(_02334_),
    .B(_02361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02404_));
 sky130_fd_sc_hd__o21a_1 _07785_ (.A1(_02365_),
    .A2(_02404_),
    .B1(_02362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02405_));
 sky130_fd_sc_hd__o21ba_1 _07786_ (.A1(_02329_),
    .A2(_02403_),
    .B1_N(_02405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02406_));
 sky130_fd_sc_hd__xor2_1 _07787_ (.A(_02401_),
    .B(_02406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02407_));
 sky130_fd_sc_hd__o22a_1 _07788_ (.A1(\sha256cu.m_out_digest.a_in[10] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(_02407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00105_));
 sky130_fd_sc_hd__or2b_1 _07789_ (.A(_02394_),
    .B_N(_02396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02408_));
 sky130_fd_sc_hd__a21boi_2 _07790_ (.A1(\sha256cu.K[10] ),
    .A2(_02397_),
    .B1_N(_02408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02409_));
 sky130_fd_sc_hd__a21o_1 _07791_ (.A1(\sha256cu.iter_processing.w[10] ),
    .A2(_02376_),
    .B1(_02375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02410_));
 sky130_fd_sc_hd__a21o_1 _07792_ (.A1(\sha256cu.m_out_digest.b_in[11] ),
    .A2(\sha256cu.m_out_digest.a_in[11] ),
    .B1(\sha256cu.m_out_digest.c_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02411_));
 sky130_fd_sc_hd__o21ai_2 _07793_ (.A1(\sha256cu.m_out_digest.b_in[11] ),
    .A2(\sha256cu.m_out_digest.a_in[11] ),
    .B1(_02411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02412_));
 sky130_fd_sc_hd__mux2_2 _07794_ (.A0(\sha256cu.m_out_digest.g_in[11] ),
    .A1(\sha256cu.m_out_digest.f_in[11] ),
    .S(\sha256cu.m_out_digest.e_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02413_));
 sky130_fd_sc_hd__xnor2_2 _07795_ (.A(_02412_),
    .B(_02413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02414_));
 sky130_fd_sc_hd__xnor2_2 _07796_ (.A(\sha256cu.iter_processing.w[11] ),
    .B(_02414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02415_));
 sky130_fd_sc_hd__xnor2_2 _07797_ (.A(\sha256cu.m_out_digest.e_in[17] ),
    .B(\sha256cu.m_out_digest.e_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02416_));
 sky130_fd_sc_hd__xnor2_2 _07798_ (.A(\sha256cu.m_out_digest.e_in[22] ),
    .B(_02416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02417_));
 sky130_fd_sc_hd__inv_2 _07799_ (.A(_02417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02418_));
 sky130_fd_sc_hd__xnor2_1 _07800_ (.A(_02027_),
    .B(\sha256cu.m_out_digest.a_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02419_));
 sky130_fd_sc_hd__xnor2_2 _07801_ (.A(_02083_),
    .B(_02419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02420_));
 sky130_fd_sc_hd__xnor2_2 _07802_ (.A(\sha256cu.m_out_digest.h_in[11] ),
    .B(_02420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02421_));
 sky130_fd_sc_hd__xnor2_2 _07803_ (.A(_02418_),
    .B(_02421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _07804_ (.A(\sha256cu.m_out_digest.h_in[10] ),
    .B(_02384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02423_));
 sky130_fd_sc_hd__o21a_1 _07805_ (.A1(_02381_),
    .A2(_02385_),
    .B1(_02423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02424_));
 sky130_fd_sc_hd__xnor2_2 _07806_ (.A(_02422_),
    .B(_02424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02425_));
 sky130_fd_sc_hd__xor2_2 _07807_ (.A(_02415_),
    .B(_02425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02426_));
 sky130_fd_sc_hd__nor2_1 _07808_ (.A(_02386_),
    .B(_02388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02427_));
 sky130_fd_sc_hd__o21ba_1 _07809_ (.A1(_02378_),
    .A2(_02389_),
    .B1_N(_02427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02428_));
 sky130_fd_sc_hd__xnor2_2 _07810_ (.A(_02426_),
    .B(_02428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02429_));
 sky130_fd_sc_hd__xnor2_2 _07811_ (.A(_02410_),
    .B(_02429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02430_));
 sky130_fd_sc_hd__and2b_1 _07812_ (.A_N(_02392_),
    .B(_02390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02431_));
 sky130_fd_sc_hd__a21oi_2 _07813_ (.A1(_02371_),
    .A2(_02393_),
    .B1(_02431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02432_));
 sky130_fd_sc_hd__xor2_2 _07814_ (.A(_02430_),
    .B(_02432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02433_));
 sky130_fd_sc_hd__xnor2_2 _07815_ (.A(\sha256cu.K[11] ),
    .B(_02433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02434_));
 sky130_fd_sc_hd__xor2_2 _07816_ (.A(_02409_),
    .B(_02434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02435_));
 sky130_fd_sc_hd__nor2_1 _07817_ (.A(_02398_),
    .B(_02400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02436_));
 sky130_fd_sc_hd__o21ba_1 _07818_ (.A1(_02401_),
    .A2(_02406_),
    .B1_N(_02436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02437_));
 sky130_fd_sc_hd__xnor2_2 _07819_ (.A(_02435_),
    .B(_02437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02438_));
 sky130_fd_sc_hd__clkbuf_4 _07820_ (.A(_02064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02439_));
 sky130_fd_sc_hd__buf_4 _07821_ (.A(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02440_));
 sky130_fd_sc_hd__or2_1 _07822_ (.A(\sha256cu.m_out_digest.a_in[11] ),
    .B(_02440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02441_));
 sky130_fd_sc_hd__o211a_1 _07823_ (.A1(_02332_),
    .A2(_02438_),
    .B1(_02441_),
    .C1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00106_));
 sky130_fd_sc_hd__and2b_1 _07824_ (.A_N(_02412_),
    .B(_02413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02442_));
 sky130_fd_sc_hd__a21o_1 _07825_ (.A1(\sha256cu.iter_processing.w[11] ),
    .A2(_02414_),
    .B1(_02442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02443_));
 sky130_fd_sc_hd__a21o_1 _07826_ (.A1(\sha256cu.m_out_digest.b_in[12] ),
    .A2(_02382_),
    .B1(\sha256cu.m_out_digest.c_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02444_));
 sky130_fd_sc_hd__o21ai_1 _07827_ (.A1(\sha256cu.m_out_digest.b_in[12] ),
    .A2(_02382_),
    .B1(_02444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02445_));
 sky130_fd_sc_hd__mux2_2 _07828_ (.A0(\sha256cu.m_out_digest.g_in[12] ),
    .A1(\sha256cu.m_out_digest.f_in[12] ),
    .S(\sha256cu.m_out_digest.e_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02446_));
 sky130_fd_sc_hd__xnor2_1 _07829_ (.A(_02445_),
    .B(_02446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02447_));
 sky130_fd_sc_hd__xnor2_1 _07830_ (.A(\sha256cu.iter_processing.w[12] ),
    .B(_02447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02448_));
 sky130_fd_sc_hd__xnor2_1 _07831_ (.A(\sha256cu.m_out_digest.e_in[18] ),
    .B(\sha256cu.m_out_digest.e_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02449_));
 sky130_fd_sc_hd__xnor2_2 _07832_ (.A(\sha256cu.m_out_digest.e_in[23] ),
    .B(_02449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02450_));
 sky130_fd_sc_hd__inv_2 _07833_ (.A(_02450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02451_));
 sky130_fd_sc_hd__xnor2_1 _07834_ (.A(\sha256cu.m_out_digest.a_in[14] ),
    .B(\sha256cu.m_out_digest.a_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02452_));
 sky130_fd_sc_hd__xnor2_2 _07835_ (.A(\sha256cu.m_out_digest.a_in[25] ),
    .B(_02452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_2 _07836_ (.A(\sha256cu.m_out_digest.h_in[12] ),
    .B(_02453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02454_));
 sky130_fd_sc_hd__xnor2_2 _07837_ (.A(_02451_),
    .B(_02454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02455_));
 sky130_fd_sc_hd__nand2_1 _07838_ (.A(\sha256cu.m_out_digest.h_in[11] ),
    .B(_02420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02456_));
 sky130_fd_sc_hd__o21a_1 _07839_ (.A1(_02418_),
    .A2(_02421_),
    .B1(_02456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02457_));
 sky130_fd_sc_hd__xnor2_1 _07840_ (.A(_02455_),
    .B(_02457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02458_));
 sky130_fd_sc_hd__xor2_1 _07841_ (.A(_02448_),
    .B(_02458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02459_));
 sky130_fd_sc_hd__nor2_1 _07842_ (.A(_02422_),
    .B(_02424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02460_));
 sky130_fd_sc_hd__o21ba_1 _07843_ (.A1(_02415_),
    .A2(_02425_),
    .B1_N(_02460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02461_));
 sky130_fd_sc_hd__xnor2_1 _07844_ (.A(_02459_),
    .B(_02461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02462_));
 sky130_fd_sc_hd__xnor2_1 _07845_ (.A(_02443_),
    .B(_02462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02463_));
 sky130_fd_sc_hd__or2b_1 _07846_ (.A(_02428_),
    .B_N(_02426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02464_));
 sky130_fd_sc_hd__a21bo_1 _07847_ (.A1(_02410_),
    .A2(_02429_),
    .B1_N(_02464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02465_));
 sky130_fd_sc_hd__xnor2_1 _07848_ (.A(_02463_),
    .B(_02465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02466_));
 sky130_fd_sc_hd__xnor2_1 _07849_ (.A(\sha256cu.K[12] ),
    .B(_02466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02467_));
 sky130_fd_sc_hd__nor2_1 _07850_ (.A(_02430_),
    .B(_02432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02468_));
 sky130_fd_sc_hd__a21o_1 _07851_ (.A1(\sha256cu.K[11] ),
    .A2(_02433_),
    .B1(_02468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02469_));
 sky130_fd_sc_hd__xor2_1 _07852_ (.A(_02467_),
    .B(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02470_));
 sky130_fd_sc_hd__and2b_1 _07853_ (.A_N(_02401_),
    .B(_02435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02471_));
 sky130_fd_sc_hd__nand2_1 _07854_ (.A(_02402_),
    .B(_02471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _07855_ (.A(_02409_),
    .B(_02434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02473_));
 sky130_fd_sc_hd__nor2_1 _07856_ (.A(_02409_),
    .B(_02434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02474_));
 sky130_fd_sc_hd__a221o_1 _07857_ (.A1(_02436_),
    .A2(_02473_),
    .B1(_02471_),
    .B2(_02405_),
    .C1(_02474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02475_));
 sky130_fd_sc_hd__o21ba_1 _07858_ (.A1(_02329_),
    .A2(_02472_),
    .B1_N(_02475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02476_));
 sky130_fd_sc_hd__nand2_1 _07859_ (.A(_02470_),
    .B(_02476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02477_));
 sky130_fd_sc_hd__buf_4 _07860_ (.A(_02108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02478_));
 sky130_fd_sc_hd__nor2_1 _07861_ (.A(_02470_),
    .B(_02476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(_02478_),
    .B(_02479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02480_));
 sky130_fd_sc_hd__a22o_1 _07863_ (.A1(_02382_),
    .A2(_02070_),
    .B1(_02477_),
    .B2(_02480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00107_));
 sky130_fd_sc_hd__and2b_1 _07864_ (.A_N(_02467_),
    .B(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02481_));
 sky130_fd_sc_hd__or2b_1 _07865_ (.A(_02463_),
    .B_N(_02465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02482_));
 sky130_fd_sc_hd__nand2_1 _07866_ (.A(\sha256cu.K[12] ),
    .B(_02466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02483_));
 sky130_fd_sc_hd__and2b_1 _07867_ (.A_N(_02445_),
    .B(_02446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02484_));
 sky130_fd_sc_hd__a21o_1 _07868_ (.A1(\sha256cu.iter_processing.w[12] ),
    .A2(_02447_),
    .B1(_02484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02485_));
 sky130_fd_sc_hd__a21o_1 _07869_ (.A1(\sha256cu.m_out_digest.b_in[13] ),
    .A2(_02027_),
    .B1(\sha256cu.m_out_digest.c_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02486_));
 sky130_fd_sc_hd__o21ai_1 _07870_ (.A1(\sha256cu.m_out_digest.b_in[13] ),
    .A2(_02027_),
    .B1(_02486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02487_));
 sky130_fd_sc_hd__mux2_2 _07871_ (.A0(\sha256cu.m_out_digest.g_in[13] ),
    .A1(\sha256cu.m_out_digest.f_in[13] ),
    .S(\sha256cu.m_out_digest.e_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02488_));
 sky130_fd_sc_hd__xnor2_1 _07872_ (.A(_02487_),
    .B(_02488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02489_));
 sky130_fd_sc_hd__xnor2_1 _07873_ (.A(\sha256cu.iter_processing.w[13] ),
    .B(_02489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02490_));
 sky130_fd_sc_hd__xnor2_2 _07874_ (.A(\sha256cu.m_out_digest.e_in[19] ),
    .B(\sha256cu.m_out_digest.e_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02491_));
 sky130_fd_sc_hd__xnor2_4 _07875_ (.A(\sha256cu.m_out_digest.e_in[24] ),
    .B(_02491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02492_));
 sky130_fd_sc_hd__inv_2 _07876_ (.A(_02492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02493_));
 sky130_fd_sc_hd__xnor2_1 _07877_ (.A(_02084_),
    .B(\sha256cu.m_out_digest.a_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02494_));
 sky130_fd_sc_hd__xnor2_2 _07878_ (.A(_02161_),
    .B(_02494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02495_));
 sky130_fd_sc_hd__xnor2_1 _07879_ (.A(\sha256cu.m_out_digest.h_in[13] ),
    .B(_02495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02496_));
 sky130_fd_sc_hd__xnor2_1 _07880_ (.A(_02493_),
    .B(_02496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02497_));
 sky130_fd_sc_hd__nand2_1 _07881_ (.A(\sha256cu.m_out_digest.h_in[12] ),
    .B(_02453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02498_));
 sky130_fd_sc_hd__o21a_1 _07882_ (.A1(_02451_),
    .A2(_02454_),
    .B1(_02498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02499_));
 sky130_fd_sc_hd__xnor2_1 _07883_ (.A(_02497_),
    .B(_02499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02500_));
 sky130_fd_sc_hd__xor2_1 _07884_ (.A(_02490_),
    .B(_02500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02501_));
 sky130_fd_sc_hd__nor2_1 _07885_ (.A(_02455_),
    .B(_02457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02502_));
 sky130_fd_sc_hd__o21ba_1 _07886_ (.A1(_02448_),
    .A2(_02458_),
    .B1_N(_02502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02503_));
 sky130_fd_sc_hd__xnor2_1 _07887_ (.A(_02501_),
    .B(_02503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02504_));
 sky130_fd_sc_hd__xnor2_1 _07888_ (.A(_02485_),
    .B(_02504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02505_));
 sky130_fd_sc_hd__and2b_1 _07889_ (.A_N(_02461_),
    .B(_02459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02506_));
 sky130_fd_sc_hd__a21oi_1 _07890_ (.A1(_02443_),
    .A2(_02462_),
    .B1(_02506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02507_));
 sky130_fd_sc_hd__xor2_1 _07891_ (.A(_02505_),
    .B(_02507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02508_));
 sky130_fd_sc_hd__xnor2_1 _07892_ (.A(\sha256cu.K[13] ),
    .B(_02508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02509_));
 sky130_fd_sc_hd__nand3_1 _07893_ (.A(_02482_),
    .B(_02483_),
    .C(_02509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02510_));
 sky130_fd_sc_hd__inv_2 _07894_ (.A(_02510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02511_));
 sky130_fd_sc_hd__a21oi_1 _07895_ (.A1(_02482_),
    .A2(_02483_),
    .B1(_02509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02512_));
 sky130_fd_sc_hd__nor2_1 _07896_ (.A(_02511_),
    .B(_02512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02513_));
 sky130_fd_sc_hd__o21ai_1 _07897_ (.A1(_02481_),
    .A2(_02479_),
    .B1(_02513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02514_));
 sky130_fd_sc_hd__buf_4 _07898_ (.A(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02515_));
 sky130_fd_sc_hd__o31a_1 _07899_ (.A1(_02481_),
    .A2(_02479_),
    .A3(_02513_),
    .B1(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02516_));
 sky130_fd_sc_hd__a221o_1 _07900_ (.A1(_02027_),
    .A2(_02220_),
    .B1(_02514_),
    .B2(_02516_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00108_));
 sky130_fd_sc_hd__and2b_1 _07901_ (.A_N(_02487_),
    .B(_02488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02517_));
 sky130_fd_sc_hd__a21o_1 _07902_ (.A1(\sha256cu.iter_processing.w[13] ),
    .A2(_02489_),
    .B1(_02517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02518_));
 sky130_fd_sc_hd__a21o_1 _07903_ (.A1(\sha256cu.m_out_digest.b_in[14] ),
    .A2(\sha256cu.m_out_digest.a_in[14] ),
    .B1(\sha256cu.m_out_digest.c_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02519_));
 sky130_fd_sc_hd__o21ai_1 _07904_ (.A1(\sha256cu.m_out_digest.b_in[14] ),
    .A2(\sha256cu.m_out_digest.a_in[14] ),
    .B1(_02519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02520_));
 sky130_fd_sc_hd__mux2_1 _07905_ (.A0(\sha256cu.m_out_digest.g_in[14] ),
    .A1(\sha256cu.m_out_digest.f_in[14] ),
    .S(\sha256cu.m_out_digest.e_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02521_));
 sky130_fd_sc_hd__xnor2_1 _07906_ (.A(_02520_),
    .B(_02521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02522_));
 sky130_fd_sc_hd__xnor2_1 _07907_ (.A(\sha256cu.iter_processing.w[14] ),
    .B(_02522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02523_));
 sky130_fd_sc_hd__xnor2_1 _07908_ (.A(\sha256cu.m_out_digest.e_in[20] ),
    .B(\sha256cu.m_out_digest.e_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02524_));
 sky130_fd_sc_hd__xnor2_2 _07909_ (.A(\sha256cu.m_out_digest.e_in[25] ),
    .B(_02524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02525_));
 sky130_fd_sc_hd__inv_2 _07910_ (.A(_02525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02526_));
 sky130_fd_sc_hd__xnor2_1 _07911_ (.A(_02128_),
    .B(\sha256cu.m_out_digest.a_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02527_));
 sky130_fd_sc_hd__xnor2_1 _07912_ (.A(\sha256cu.m_out_digest.a_in[27] ),
    .B(_02527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02528_));
 sky130_fd_sc_hd__xnor2_1 _07913_ (.A(\sha256cu.m_out_digest.h_in[14] ),
    .B(_02528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02529_));
 sky130_fd_sc_hd__xnor2_1 _07914_ (.A(_02526_),
    .B(_02529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02530_));
 sky130_fd_sc_hd__nand2_1 _07915_ (.A(\sha256cu.m_out_digest.h_in[13] ),
    .B(_02495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02531_));
 sky130_fd_sc_hd__o21a_1 _07916_ (.A1(_02493_),
    .A2(_02496_),
    .B1(_02531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02532_));
 sky130_fd_sc_hd__xnor2_1 _07917_ (.A(_02530_),
    .B(_02532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02533_));
 sky130_fd_sc_hd__xor2_1 _07918_ (.A(_02523_),
    .B(_02533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02534_));
 sky130_fd_sc_hd__nor2_1 _07919_ (.A(_02497_),
    .B(_02499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02535_));
 sky130_fd_sc_hd__o21ba_1 _07920_ (.A1(_02490_),
    .A2(_02500_),
    .B1_N(_02535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02536_));
 sky130_fd_sc_hd__xnor2_1 _07921_ (.A(_02534_),
    .B(_02536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02537_));
 sky130_fd_sc_hd__xnor2_1 _07922_ (.A(_02518_),
    .B(_02537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02538_));
 sky130_fd_sc_hd__or2b_1 _07923_ (.A(_02503_),
    .B_N(_02501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02539_));
 sky130_fd_sc_hd__a21bo_1 _07924_ (.A1(_02485_),
    .A2(_02504_),
    .B1_N(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02540_));
 sky130_fd_sc_hd__xnor2_1 _07925_ (.A(_02538_),
    .B(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02541_));
 sky130_fd_sc_hd__xnor2_2 _07926_ (.A(\sha256cu.K[14] ),
    .B(_02541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_1 _07927_ (.A(_02505_),
    .B(_02507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02543_));
 sky130_fd_sc_hd__a21o_1 _07928_ (.A1(\sha256cu.K[13] ),
    .A2(_02508_),
    .B1(_02543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02544_));
 sky130_fd_sc_hd__xor2_2 _07929_ (.A(_02542_),
    .B(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02545_));
 sky130_fd_sc_hd__nor3b_1 _07930_ (.A(_02512_),
    .B(_02470_),
    .C_N(_02510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02546_));
 sky130_fd_sc_hd__inv_2 _07931_ (.A(_02546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02547_));
 sky130_fd_sc_hd__o21a_1 _07932_ (.A1(_02481_),
    .A2(_02512_),
    .B1(_02510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02548_));
 sky130_fd_sc_hd__o21bai_1 _07933_ (.A1(_02476_),
    .A2(_02547_),
    .B1_N(_02548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02549_));
 sky130_fd_sc_hd__xnor2_1 _07934_ (.A(_02545_),
    .B(_02549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02550_));
 sky130_fd_sc_hd__a22o_1 _07935_ (.A1(\sha256cu.m_out_digest.a_in[14] ),
    .A2(_02037_),
    .B1(_02017_),
    .B2(_02550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02551_));
 sky130_fd_sc_hd__or2_1 _07936_ (.A(_02002_),
    .B(_02551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02552_));
 sky130_fd_sc_hd__clkbuf_1 _07937_ (.A(_02552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00109_));
 sky130_fd_sc_hd__and2b_1 _07938_ (.A_N(_02542_),
    .B(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02553_));
 sky130_fd_sc_hd__and2b_1 _07939_ (.A_N(_02545_),
    .B(_02549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02554_));
 sky130_fd_sc_hd__or2b_1 _07940_ (.A(_02538_),
    .B_N(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _07941_ (.A(\sha256cu.K[14] ),
    .B(_02541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02556_));
 sky130_fd_sc_hd__and2b_1 _07942_ (.A_N(_02520_),
    .B(_02521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02557_));
 sky130_fd_sc_hd__a21o_1 _07943_ (.A1(\sha256cu.iter_processing.w[14] ),
    .A2(_02522_),
    .B1(_02557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02558_));
 sky130_fd_sc_hd__a21o_1 _07944_ (.A1(\sha256cu.m_out_digest.b_in[15] ),
    .A2(_02084_),
    .B1(\sha256cu.m_out_digest.c_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02559_));
 sky130_fd_sc_hd__o21ai_2 _07945_ (.A1(\sha256cu.m_out_digest.b_in[15] ),
    .A2(_02084_),
    .B1(_02559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02560_));
 sky130_fd_sc_hd__mux2_2 _07946_ (.A0(\sha256cu.m_out_digest.g_in[15] ),
    .A1(\sha256cu.m_out_digest.f_in[15] ),
    .S(\sha256cu.m_out_digest.e_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02561_));
 sky130_fd_sc_hd__xnor2_2 _07947_ (.A(_02560_),
    .B(_02561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02562_));
 sky130_fd_sc_hd__xnor2_2 _07948_ (.A(\sha256cu.iter_processing.w[15] ),
    .B(_02562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02563_));
 sky130_fd_sc_hd__xnor2_1 _07949_ (.A(\sha256cu.m_out_digest.e_in[21] ),
    .B(\sha256cu.m_out_digest.e_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02564_));
 sky130_fd_sc_hd__xnor2_2 _07950_ (.A(\sha256cu.m_out_digest.e_in[26] ),
    .B(_02564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02565_));
 sky130_fd_sc_hd__inv_2 _07951_ (.A(_02565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02566_));
 sky130_fd_sc_hd__xnor2_1 _07952_ (.A(_02162_),
    .B(\sha256cu.m_out_digest.a_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02567_));
 sky130_fd_sc_hd__xnor2_2 _07953_ (.A(_02232_),
    .B(_02567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02568_));
 sky130_fd_sc_hd__xnor2_2 _07954_ (.A(\sha256cu.m_out_digest.h_in[15] ),
    .B(_02568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02569_));
 sky130_fd_sc_hd__xnor2_2 _07955_ (.A(_02566_),
    .B(_02569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _07956_ (.A(\sha256cu.m_out_digest.h_in[14] ),
    .B(_02528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02571_));
 sky130_fd_sc_hd__o21a_1 _07957_ (.A1(_02526_),
    .A2(_02529_),
    .B1(_02571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02572_));
 sky130_fd_sc_hd__xnor2_2 _07958_ (.A(_02570_),
    .B(_02572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02573_));
 sky130_fd_sc_hd__xor2_2 _07959_ (.A(_02563_),
    .B(_02573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02574_));
 sky130_fd_sc_hd__nor2_1 _07960_ (.A(_02530_),
    .B(_02532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02575_));
 sky130_fd_sc_hd__o21bai_2 _07961_ (.A1(_02523_),
    .A2(_02533_),
    .B1_N(_02575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02576_));
 sky130_fd_sc_hd__xor2_2 _07962_ (.A(_02574_),
    .B(_02576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02577_));
 sky130_fd_sc_hd__xnor2_2 _07963_ (.A(_02558_),
    .B(_02577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02578_));
 sky130_fd_sc_hd__and2b_1 _07964_ (.A_N(_02536_),
    .B(_02534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02579_));
 sky130_fd_sc_hd__a21oi_2 _07965_ (.A1(_02518_),
    .A2(_02537_),
    .B1(_02579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02580_));
 sky130_fd_sc_hd__xor2_2 _07966_ (.A(_02578_),
    .B(_02580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02581_));
 sky130_fd_sc_hd__xnor2_2 _07967_ (.A(\sha256cu.K[15] ),
    .B(_02581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02582_));
 sky130_fd_sc_hd__nand3_2 _07968_ (.A(_02555_),
    .B(_02556_),
    .C(_02582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02583_));
 sky130_fd_sc_hd__inv_2 _07969_ (.A(_02583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02584_));
 sky130_fd_sc_hd__a21oi_2 _07970_ (.A1(_02555_),
    .A2(_02556_),
    .B1(_02582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02585_));
 sky130_fd_sc_hd__nor2_1 _07971_ (.A(_02584_),
    .B(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02586_));
 sky130_fd_sc_hd__o21ai_1 _07972_ (.A1(_02553_),
    .A2(_02554_),
    .B1(_02586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02587_));
 sky130_fd_sc_hd__o31a_1 _07973_ (.A1(_02553_),
    .A2(_02554_),
    .A3(_02586_),
    .B1(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02588_));
 sky130_fd_sc_hd__a221o_1 _07974_ (.A1(_02084_),
    .A2(_02220_),
    .B1(_02587_),
    .B2(_02588_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00110_));
 sky130_fd_sc_hd__or2_1 _07975_ (.A(_02578_),
    .B(_02580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02589_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(\sha256cu.K[15] ),
    .B(_02581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02590_));
 sky130_fd_sc_hd__and2b_1 _07977_ (.A_N(_02560_),
    .B(_02561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02591_));
 sky130_fd_sc_hd__a21o_1 _07978_ (.A1(\sha256cu.iter_processing.w[15] ),
    .A2(_02562_),
    .B1(_02591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02592_));
 sky130_fd_sc_hd__a21o_1 _07979_ (.A1(\sha256cu.m_out_digest.b_in[16] ),
    .A2(_02128_),
    .B1(\sha256cu.m_out_digest.c_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02593_));
 sky130_fd_sc_hd__o21ai_1 _07980_ (.A1(\sha256cu.m_out_digest.b_in[16] ),
    .A2(_02128_),
    .B1(_02593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02594_));
 sky130_fd_sc_hd__mux2_2 _07981_ (.A0(\sha256cu.m_out_digest.g_in[16] ),
    .A1(\sha256cu.m_out_digest.f_in[16] ),
    .S(\sha256cu.m_out_digest.e_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02595_));
 sky130_fd_sc_hd__xnor2_1 _07982_ (.A(_02594_),
    .B(_02595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02596_));
 sky130_fd_sc_hd__xnor2_1 _07983_ (.A(\sha256cu.iter_processing.w[16] ),
    .B(_02596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02597_));
 sky130_fd_sc_hd__xnor2_1 _07984_ (.A(\sha256cu.m_out_digest.e_in[22] ),
    .B(\sha256cu.m_out_digest.e_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02598_));
 sky130_fd_sc_hd__xnor2_2 _07985_ (.A(\sha256cu.m_out_digest.e_in[27] ),
    .B(_02598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02599_));
 sky130_fd_sc_hd__inv_2 _07986_ (.A(_02599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02600_));
 sky130_fd_sc_hd__xnor2_1 _07987_ (.A(_02198_),
    .B(\sha256cu.m_out_digest.a_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02601_));
 sky130_fd_sc_hd__xnor2_2 _07988_ (.A(_02272_),
    .B(_02601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02602_));
 sky130_fd_sc_hd__xnor2_1 _07989_ (.A(\sha256cu.m_out_digest.h_in[16] ),
    .B(_02602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02603_));
 sky130_fd_sc_hd__xnor2_1 _07990_ (.A(_02600_),
    .B(_02603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02604_));
 sky130_fd_sc_hd__nand2_1 _07991_ (.A(\sha256cu.m_out_digest.h_in[15] ),
    .B(_02568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02605_));
 sky130_fd_sc_hd__o21a_1 _07992_ (.A1(_02566_),
    .A2(_02569_),
    .B1(_02605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02606_));
 sky130_fd_sc_hd__xnor2_1 _07993_ (.A(_02604_),
    .B(_02606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02607_));
 sky130_fd_sc_hd__xor2_1 _07994_ (.A(_02597_),
    .B(_02607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02608_));
 sky130_fd_sc_hd__nor2_1 _07995_ (.A(_02570_),
    .B(_02572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02609_));
 sky130_fd_sc_hd__o21ba_1 _07996_ (.A1(_02563_),
    .A2(_02573_),
    .B1_N(_02609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02610_));
 sky130_fd_sc_hd__xnor2_1 _07997_ (.A(_02608_),
    .B(_02610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02611_));
 sky130_fd_sc_hd__xnor2_1 _07998_ (.A(_02592_),
    .B(_02611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02612_));
 sky130_fd_sc_hd__and2_1 _07999_ (.A(_02574_),
    .B(_02576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02613_));
 sky130_fd_sc_hd__a21o_1 _08000_ (.A1(_02558_),
    .A2(_02577_),
    .B1(_02613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02614_));
 sky130_fd_sc_hd__xnor2_1 _08001_ (.A(_02612_),
    .B(_02614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02615_));
 sky130_fd_sc_hd__or2_1 _08002_ (.A(\sha256cu.K[16] ),
    .B(_02615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02616_));
 sky130_fd_sc_hd__nand2_1 _08003_ (.A(\sha256cu.K[16] ),
    .B(_02615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02617_));
 sky130_fd_sc_hd__nand2_1 _08004_ (.A(_02616_),
    .B(_02617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02618_));
 sky130_fd_sc_hd__a21oi_2 _08005_ (.A1(_02589_),
    .A2(_02590_),
    .B1(_02618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02619_));
 sky130_fd_sc_hd__and3_1 _08006_ (.A(_02589_),
    .B(_02590_),
    .C(_02618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02620_));
 sky130_fd_sc_hd__or2_1 _08007_ (.A(_02619_),
    .B(_02620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02621_));
 sky130_fd_sc_hd__nor3b_2 _08008_ (.A(_02585_),
    .B(_02545_),
    .C_N(_02583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02622_));
 sky130_fd_sc_hd__a221oi_4 _08009_ (.A1(_02553_),
    .A2(_02583_),
    .B1(_02622_),
    .B2(_02548_),
    .C1(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02623_));
 sky130_fd_sc_hd__and2_1 _08010_ (.A(_02546_),
    .B(_02622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02624_));
 sky130_fd_sc_hd__nand4_1 _08011_ (.A(_02402_),
    .B(_02471_),
    .C(_02546_),
    .D(_02622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02625_));
 sky130_fd_sc_hd__o2bb2a_1 _08012_ (.A1_N(_02475_),
    .A2_N(_02624_),
    .B1(_02625_),
    .B2(_02329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02626_));
 sky130_fd_sc_hd__and2_1 _08013_ (.A(_02623_),
    .B(_02626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02627_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(_02621_),
    .B(_02627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02628_));
 sky130_fd_sc_hd__buf_4 _08015_ (.A(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02629_));
 sky130_fd_sc_hd__nor2_2 _08016_ (.A(_02621_),
    .B(_02627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02630_));
 sky130_fd_sc_hd__nor2_1 _08017_ (.A(_02629_),
    .B(_02630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02631_));
 sky130_fd_sc_hd__a221o_1 _08018_ (.A1(_02128_),
    .A2(_02220_),
    .B1(_02628_),
    .B2(_02631_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00111_));
 sky130_fd_sc_hd__or2b_1 _08019_ (.A(_02612_),
    .B_N(_02614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02632_));
 sky130_fd_sc_hd__or2b_1 _08020_ (.A(_02610_),
    .B_N(_02608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02633_));
 sky130_fd_sc_hd__a21bo_1 _08021_ (.A1(_02592_),
    .A2(_02611_),
    .B1_N(_02633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02634_));
 sky130_fd_sc_hd__and2b_1 _08022_ (.A_N(_02594_),
    .B(_02595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02635_));
 sky130_fd_sc_hd__a21o_1 _08023_ (.A1(\sha256cu.iter_processing.w[16] ),
    .A2(_02596_),
    .B1(_02635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02636_));
 sky130_fd_sc_hd__a21o_1 _08024_ (.A1(\sha256cu.m_out_digest.b_in[17] ),
    .A2(_02162_),
    .B1(\sha256cu.m_out_digest.c_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02637_));
 sky130_fd_sc_hd__o21ai_1 _08025_ (.A1(\sha256cu.m_out_digest.b_in[17] ),
    .A2(_02162_),
    .B1(_02637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02638_));
 sky130_fd_sc_hd__mux2_1 _08026_ (.A0(\sha256cu.m_out_digest.g_in[17] ),
    .A1(\sha256cu.m_out_digest.f_in[17] ),
    .S(\sha256cu.m_out_digest.e_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02639_));
 sky130_fd_sc_hd__xnor2_1 _08027_ (.A(_02638_),
    .B(_02639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02640_));
 sky130_fd_sc_hd__xnor2_1 _08028_ (.A(\sha256cu.iter_processing.w[17] ),
    .B(_02640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02641_));
 sky130_fd_sc_hd__xnor2_2 _08029_ (.A(\sha256cu.m_out_digest.e_in[23] ),
    .B(\sha256cu.m_out_digest.e_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02642_));
 sky130_fd_sc_hd__xnor2_4 _08030_ (.A(\sha256cu.m_out_digest.e_in[28] ),
    .B(_02642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02643_));
 sky130_fd_sc_hd__inv_2 _08031_ (.A(_02643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02644_));
 sky130_fd_sc_hd__xnor2_1 _08032_ (.A(_02233_),
    .B(\sha256cu.m_out_digest.a_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02645_));
 sky130_fd_sc_hd__xnor2_2 _08033_ (.A(_02304_),
    .B(_02645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02646_));
 sky130_fd_sc_hd__xnor2_1 _08034_ (.A(\sha256cu.m_out_digest.h_in[17] ),
    .B(_02646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02647_));
 sky130_fd_sc_hd__xnor2_1 _08035_ (.A(_02644_),
    .B(_02647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02648_));
 sky130_fd_sc_hd__nand2_1 _08036_ (.A(\sha256cu.m_out_digest.h_in[16] ),
    .B(_02602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02649_));
 sky130_fd_sc_hd__o21a_1 _08037_ (.A1(_02600_),
    .A2(_02603_),
    .B1(_02649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02650_));
 sky130_fd_sc_hd__xnor2_1 _08038_ (.A(_02648_),
    .B(_02650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02651_));
 sky130_fd_sc_hd__xor2_1 _08039_ (.A(_02641_),
    .B(_02651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02652_));
 sky130_fd_sc_hd__or2_1 _08040_ (.A(_02597_),
    .B(_02607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02653_));
 sky130_fd_sc_hd__o21a_1 _08041_ (.A1(_02604_),
    .A2(_02606_),
    .B1(_02653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02654_));
 sky130_fd_sc_hd__xnor2_1 _08042_ (.A(_02652_),
    .B(_02654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02655_));
 sky130_fd_sc_hd__xnor2_1 _08043_ (.A(_02636_),
    .B(_02655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02656_));
 sky130_fd_sc_hd__xnor2_1 _08044_ (.A(_02634_),
    .B(_02656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02657_));
 sky130_fd_sc_hd__xnor2_1 _08045_ (.A(\sha256cu.K[17] ),
    .B(_02657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02658_));
 sky130_fd_sc_hd__and3_1 _08046_ (.A(_02632_),
    .B(_02617_),
    .C(_02658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02659_));
 sky130_fd_sc_hd__a21oi_1 _08047_ (.A1(_02632_),
    .A2(_02617_),
    .B1(_02658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02660_));
 sky130_fd_sc_hd__or2_2 _08048_ (.A(_02659_),
    .B(_02660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02661_));
 sky130_fd_sc_hd__o21ai_1 _08049_ (.A1(_02619_),
    .A2(_02630_),
    .B1(_02661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02662_));
 sky130_fd_sc_hd__o31a_1 _08050_ (.A1(_02619_),
    .A2(_02630_),
    .A3(_02661_),
    .B1(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02663_));
 sky130_fd_sc_hd__o21ai_1 _08051_ (.A1(_02162_),
    .A2(_02440_),
    .B1(_01966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02664_));
 sky130_fd_sc_hd__a21oi_1 _08052_ (.A1(_02662_),
    .A2(_02663_),
    .B1(_02664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00112_));
 sky130_fd_sc_hd__or2b_1 _08053_ (.A(_02654_),
    .B_N(_02652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02665_));
 sky130_fd_sc_hd__a21bo_1 _08054_ (.A1(_02636_),
    .A2(_02655_),
    .B1_N(_02665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02666_));
 sky130_fd_sc_hd__and2b_1 _08055_ (.A_N(_02638_),
    .B(_02639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02667_));
 sky130_fd_sc_hd__a21o_1 _08056_ (.A1(\sha256cu.iter_processing.w[17] ),
    .A2(_02640_),
    .B1(_02667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02668_));
 sky130_fd_sc_hd__a21o_1 _08057_ (.A1(\sha256cu.m_out_digest.b_in[18] ),
    .A2(_02198_),
    .B1(\sha256cu.m_out_digest.c_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02669_));
 sky130_fd_sc_hd__o21ai_1 _08058_ (.A1(\sha256cu.m_out_digest.b_in[18] ),
    .A2(_02198_),
    .B1(_02669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02670_));
 sky130_fd_sc_hd__mux2_1 _08059_ (.A0(\sha256cu.m_out_digest.g_in[18] ),
    .A1(\sha256cu.m_out_digest.f_in[18] ),
    .S(\sha256cu.m_out_digest.e_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02671_));
 sky130_fd_sc_hd__xnor2_1 _08060_ (.A(_02670_),
    .B(_02671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02672_));
 sky130_fd_sc_hd__xnor2_1 _08061_ (.A(\sha256cu.iter_processing.w[18] ),
    .B(_02672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02673_));
 sky130_fd_sc_hd__xnor2_2 _08062_ (.A(\sha256cu.m_out_digest.e_in[24] ),
    .B(\sha256cu.m_out_digest.e_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02674_));
 sky130_fd_sc_hd__xnor2_4 _08063_ (.A(\sha256cu.m_out_digest.e_in[29] ),
    .B(_02674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02675_));
 sky130_fd_sc_hd__inv_2 _08064_ (.A(_02675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02676_));
 sky130_fd_sc_hd__xnor2_1 _08065_ (.A(_02273_),
    .B(\sha256cu.m_out_digest.a_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02677_));
 sky130_fd_sc_hd__xnor2_2 _08066_ (.A(\sha256cu.m_out_digest.a_in[31] ),
    .B(_02677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02678_));
 sky130_fd_sc_hd__xnor2_1 _08067_ (.A(\sha256cu.m_out_digest.h_in[18] ),
    .B(_02678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02679_));
 sky130_fd_sc_hd__xnor2_1 _08068_ (.A(_02676_),
    .B(_02679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02680_));
 sky130_fd_sc_hd__nand2_1 _08069_ (.A(\sha256cu.m_out_digest.h_in[17] ),
    .B(_02646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02681_));
 sky130_fd_sc_hd__o21a_1 _08070_ (.A1(_02644_),
    .A2(_02647_),
    .B1(_02681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02682_));
 sky130_fd_sc_hd__xnor2_1 _08071_ (.A(_02680_),
    .B(_02682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02683_));
 sky130_fd_sc_hd__xor2_1 _08072_ (.A(_02673_),
    .B(_02683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02684_));
 sky130_fd_sc_hd__nor2_1 _08073_ (.A(_02648_),
    .B(_02650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02685_));
 sky130_fd_sc_hd__o21bai_2 _08074_ (.A1(_02641_),
    .A2(_02651_),
    .B1_N(_02685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02686_));
 sky130_fd_sc_hd__xor2_1 _08075_ (.A(_02684_),
    .B(_02686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02687_));
 sky130_fd_sc_hd__and2_1 _08076_ (.A(_02668_),
    .B(_02687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02688_));
 sky130_fd_sc_hd__nor2_1 _08077_ (.A(_02668_),
    .B(_02687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02689_));
 sky130_fd_sc_hd__or2_1 _08078_ (.A(_02688_),
    .B(_02689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02690_));
 sky130_fd_sc_hd__xnor2_2 _08079_ (.A(_02666_),
    .B(_02690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02691_));
 sky130_fd_sc_hd__xnor2_2 _08080_ (.A(\sha256cu.K[18] ),
    .B(_02691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02692_));
 sky130_fd_sc_hd__or2b_1 _08081_ (.A(_02656_),
    .B_N(_02634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02693_));
 sky130_fd_sc_hd__a21bo_1 _08082_ (.A1(\sha256cu.K[17] ),
    .A2(_02657_),
    .B1_N(_02693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02694_));
 sky130_fd_sc_hd__xor2_2 _08083_ (.A(_02692_),
    .B(_02694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02695_));
 sky130_fd_sc_hd__inv_2 _08084_ (.A(_02661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02696_));
 sky130_fd_sc_hd__o21ba_1 _08085_ (.A1(_02619_),
    .A2(_02660_),
    .B1_N(_02659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02697_));
 sky130_fd_sc_hd__a21oi_2 _08086_ (.A1(_02630_),
    .A2(_02696_),
    .B1(_02697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02698_));
 sky130_fd_sc_hd__a21oi_1 _08087_ (.A1(_02695_),
    .A2(_02698_),
    .B1(_02108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02699_));
 sky130_fd_sc_hd__o21a_1 _08088_ (.A1(_02695_),
    .A2(_02698_),
    .B1(_02699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02700_));
 sky130_fd_sc_hd__a21o_1 _08089_ (.A1(_02198_),
    .A2(_02070_),
    .B1(_02700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00113_));
 sky130_fd_sc_hd__or2b_1 _08090_ (.A(_02690_),
    .B_N(_02666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02701_));
 sky130_fd_sc_hd__a21boi_2 _08091_ (.A1(\sha256cu.K[18] ),
    .A2(_02691_),
    .B1_N(_02701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02702_));
 sky130_fd_sc_hd__a21oi_2 _08092_ (.A1(_02684_),
    .A2(_02686_),
    .B1(_02688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02703_));
 sky130_fd_sc_hd__and2b_1 _08093_ (.A_N(_02670_),
    .B(_02671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02704_));
 sky130_fd_sc_hd__a21o_1 _08094_ (.A1(\sha256cu.iter_processing.w[18] ),
    .A2(_02672_),
    .B1(_02704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02705_));
 sky130_fd_sc_hd__a21o_1 _08095_ (.A1(\sha256cu.m_out_digest.b_in[19] ),
    .A2(_02233_),
    .B1(\sha256cu.m_out_digest.c_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02706_));
 sky130_fd_sc_hd__o21ai_2 _08096_ (.A1(\sha256cu.m_out_digest.b_in[19] ),
    .A2(_02233_),
    .B1(_02706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02707_));
 sky130_fd_sc_hd__mux2_2 _08097_ (.A0(\sha256cu.m_out_digest.g_in[19] ),
    .A1(\sha256cu.m_out_digest.f_in[19] ),
    .S(\sha256cu.m_out_digest.e_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02708_));
 sky130_fd_sc_hd__xnor2_1 _08098_ (.A(_02707_),
    .B(_02708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02709_));
 sky130_fd_sc_hd__xnor2_1 _08099_ (.A(\sha256cu.iter_processing.w[19] ),
    .B(_02709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02710_));
 sky130_fd_sc_hd__xnor2_2 _08100_ (.A(\sha256cu.m_out_digest.e_in[25] ),
    .B(\sha256cu.m_out_digest.e_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02711_));
 sky130_fd_sc_hd__xnor2_2 _08101_ (.A(\sha256cu.m_out_digest.e_in[30] ),
    .B(_02711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02712_));
 sky130_fd_sc_hd__inv_2 _08102_ (.A(_02712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02713_));
 sky130_fd_sc_hd__xnor2_1 _08103_ (.A(\sha256cu.m_out_digest.a_in[9] ),
    .B(\sha256cu.m_out_digest.a_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02714_));
 sky130_fd_sc_hd__xnor2_1 _08104_ (.A(\sha256cu.m_out_digest.a_in[21] ),
    .B(_02714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02715_));
 sky130_fd_sc_hd__xnor2_1 _08105_ (.A(\sha256cu.m_out_digest.h_in[19] ),
    .B(_02715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02716_));
 sky130_fd_sc_hd__xnor2_1 _08106_ (.A(_02713_),
    .B(_02716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02717_));
 sky130_fd_sc_hd__nand2_1 _08107_ (.A(\sha256cu.m_out_digest.h_in[18] ),
    .B(_02678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02718_));
 sky130_fd_sc_hd__o21a_1 _08108_ (.A1(_02676_),
    .A2(_02679_),
    .B1(_02718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02719_));
 sky130_fd_sc_hd__xnor2_1 _08109_ (.A(_02717_),
    .B(_02719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02720_));
 sky130_fd_sc_hd__xor2_1 _08110_ (.A(_02710_),
    .B(_02720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02721_));
 sky130_fd_sc_hd__or2_1 _08111_ (.A(_02673_),
    .B(_02683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02722_));
 sky130_fd_sc_hd__o21a_1 _08112_ (.A1(_02680_),
    .A2(_02682_),
    .B1(_02722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02723_));
 sky130_fd_sc_hd__xnor2_1 _08113_ (.A(_02721_),
    .B(_02723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02724_));
 sky130_fd_sc_hd__xnor2_1 _08114_ (.A(_02705_),
    .B(_02724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02725_));
 sky130_fd_sc_hd__xor2_2 _08115_ (.A(_02703_),
    .B(_02725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02726_));
 sky130_fd_sc_hd__xnor2_2 _08116_ (.A(\sha256cu.K[19] ),
    .B(_02726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02727_));
 sky130_fd_sc_hd__xor2_1 _08117_ (.A(_02702_),
    .B(_02727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02728_));
 sky130_fd_sc_hd__and2b_1 _08118_ (.A_N(_02692_),
    .B(_02694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02729_));
 sky130_fd_sc_hd__o21ba_1 _08119_ (.A1(_02695_),
    .A2(_02698_),
    .B1_N(_02729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02730_));
 sky130_fd_sc_hd__xor2_1 _08120_ (.A(_02728_),
    .B(_02730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02731_));
 sky130_fd_sc_hd__buf_4 _08121_ (.A(_02037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02732_));
 sky130_fd_sc_hd__nand2_1 _08122_ (.A(_02233_),
    .B(_02732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02733_));
 sky130_fd_sc_hd__o211ai_1 _08123_ (.A1(_02332_),
    .A2(_02731_),
    .B1(_02733_),
    .C1(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00114_));
 sky130_fd_sc_hd__or2b_1 _08124_ (.A(_02723_),
    .B_N(_02721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02734_));
 sky130_fd_sc_hd__a21bo_1 _08125_ (.A1(_02705_),
    .A2(_02724_),
    .B1_N(_02734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02735_));
 sky130_fd_sc_hd__and2b_1 _08126_ (.A_N(_02707_),
    .B(_02708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02736_));
 sky130_fd_sc_hd__a21o_1 _08127_ (.A1(\sha256cu.iter_processing.w[19] ),
    .A2(_02709_),
    .B1(_02736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02737_));
 sky130_fd_sc_hd__a21o_1 _08128_ (.A1(\sha256cu.m_out_digest.b_in[20] ),
    .A2(_02273_),
    .B1(\sha256cu.m_out_digest.c_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02738_));
 sky130_fd_sc_hd__o21ai_2 _08129_ (.A1(\sha256cu.m_out_digest.b_in[20] ),
    .A2(_02273_),
    .B1(_02738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02739_));
 sky130_fd_sc_hd__mux2_2 _08130_ (.A0(\sha256cu.m_out_digest.g_in[20] ),
    .A1(\sha256cu.m_out_digest.f_in[20] ),
    .S(\sha256cu.m_out_digest.e_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02740_));
 sky130_fd_sc_hd__xnor2_2 _08131_ (.A(_02739_),
    .B(_02740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02741_));
 sky130_fd_sc_hd__xor2_2 _08132_ (.A(\sha256cu.iter_processing.w[20] ),
    .B(_02741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02742_));
 sky130_fd_sc_hd__xnor2_2 _08133_ (.A(\sha256cu.m_out_digest.a_in[10] ),
    .B(\sha256cu.m_out_digest.a_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02743_));
 sky130_fd_sc_hd__xnor2_2 _08134_ (.A(_02026_),
    .B(_02743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02744_));
 sky130_fd_sc_hd__xnor2_2 _08135_ (.A(\sha256cu.m_out_digest.h_in[20] ),
    .B(_02744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02745_));
 sky130_fd_sc_hd__xnor2_2 _08136_ (.A(\sha256cu.m_out_digest.e_in[26] ),
    .B(\sha256cu.m_out_digest.e_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor2_4 _08137_ (.A(\sha256cu.m_out_digest.e_in[31] ),
    .B(_02746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02747_));
 sky130_fd_sc_hd__xnor2_2 _08138_ (.A(_02745_),
    .B(_02747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02748_));
 sky130_fd_sc_hd__nand2_1 _08139_ (.A(\sha256cu.m_out_digest.h_in[19] ),
    .B(_02715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02749_));
 sky130_fd_sc_hd__o21a_1 _08140_ (.A1(_02713_),
    .A2(_02716_),
    .B1(_02749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02750_));
 sky130_fd_sc_hd__xnor2_2 _08141_ (.A(_02748_),
    .B(_02750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02751_));
 sky130_fd_sc_hd__xor2_2 _08142_ (.A(_02742_),
    .B(_02751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02752_));
 sky130_fd_sc_hd__nor2_1 _08143_ (.A(_02717_),
    .B(_02719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02753_));
 sky130_fd_sc_hd__o21ba_1 _08144_ (.A1(_02710_),
    .A2(_02720_),
    .B1_N(_02753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02754_));
 sky130_fd_sc_hd__xnor2_2 _08145_ (.A(_02752_),
    .B(_02754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02755_));
 sky130_fd_sc_hd__xnor2_2 _08146_ (.A(_02737_),
    .B(_02755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_2 _08147_ (.A(_02735_),
    .B(_02756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02757_));
 sky130_fd_sc_hd__xnor2_2 _08148_ (.A(\sha256cu.K[20] ),
    .B(_02757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02758_));
 sky130_fd_sc_hd__nor2_1 _08149_ (.A(_02703_),
    .B(_02725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02759_));
 sky130_fd_sc_hd__a21oi_2 _08150_ (.A1(\sha256cu.K[19] ),
    .A2(_02726_),
    .B1(_02759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02760_));
 sky130_fd_sc_hd__xnor2_2 _08151_ (.A(_02758_),
    .B(_02760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02761_));
 sky130_fd_sc_hd__and2b_1 _08152_ (.A_N(_02695_),
    .B(_02728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02762_));
 sky130_fd_sc_hd__or3b_1 _08153_ (.A(_02621_),
    .B(_02661_),
    .C_N(_02762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02763_));
 sky130_fd_sc_hd__nand2_1 _08154_ (.A(_02702_),
    .B(_02727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02764_));
 sky130_fd_sc_hd__nor2_1 _08155_ (.A(_02702_),
    .B(_02727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02765_));
 sky130_fd_sc_hd__a221oi_4 _08156_ (.A1(_02729_),
    .A2(_02764_),
    .B1(_02762_),
    .B2(_02697_),
    .C1(_02765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02766_));
 sky130_fd_sc_hd__o21a_1 _08157_ (.A1(_02627_),
    .A2(_02763_),
    .B1(_02766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_1 _08158_ (.A(_02761_),
    .B(_02767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02768_));
 sky130_fd_sc_hd__a21o_1 _08159_ (.A1(_02761_),
    .A2(_02767_),
    .B1(_02478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02769_));
 sky130_fd_sc_hd__a2bb2o_1 _08160_ (.A1_N(_02768_),
    .A2_N(_02769_),
    .B1(_02273_),
    .B2(_02070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00115_));
 sky130_fd_sc_hd__and2b_1 _08161_ (.A_N(_02739_),
    .B(_02740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02770_));
 sky130_fd_sc_hd__a21o_1 _08162_ (.A1(\sha256cu.iter_processing.w[20] ),
    .A2(_02741_),
    .B1(_02770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02771_));
 sky130_fd_sc_hd__inv_2 _08163_ (.A(_02771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02772_));
 sky130_fd_sc_hd__xnor2_2 _08164_ (.A(\sha256cu.m_out_digest.a_in[11] ),
    .B(\sha256cu.m_out_digest.a_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02773_));
 sky130_fd_sc_hd__xnor2_1 _08165_ (.A(\sha256cu.m_out_digest.a_in[23] ),
    .B(_02773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02774_));
 sky130_fd_sc_hd__xnor2_1 _08166_ (.A(\sha256cu.m_out_digest.h_in[21] ),
    .B(_02774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02775_));
 sky130_fd_sc_hd__xnor2_4 _08167_ (.A(\sha256cu.m_out_digest.e_in[14] ),
    .B(\sha256cu.m_out_digest.e_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02776_));
 sky130_fd_sc_hd__xnor2_4 _08168_ (.A(\sha256cu.m_out_digest.e_in[27] ),
    .B(_02776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02777_));
 sky130_fd_sc_hd__xnor2_1 _08169_ (.A(_02775_),
    .B(_02777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02778_));
 sky130_fd_sc_hd__inv_2 _08170_ (.A(_02747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02779_));
 sky130_fd_sc_hd__nand2_1 _08171_ (.A(\sha256cu.m_out_digest.h_in[20] ),
    .B(_02744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02780_));
 sky130_fd_sc_hd__o21ai_1 _08172_ (.A1(_02745_),
    .A2(_02779_),
    .B1(_02780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02781_));
 sky130_fd_sc_hd__xor2_1 _08173_ (.A(_02778_),
    .B(_02781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02782_));
 sky130_fd_sc_hd__a21o_1 _08174_ (.A1(\sha256cu.m_out_digest.b_in[21] ),
    .A2(\sha256cu.m_out_digest.a_in[21] ),
    .B1(\sha256cu.m_out_digest.c_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02783_));
 sky130_fd_sc_hd__o21ai_1 _08175_ (.A1(\sha256cu.m_out_digest.b_in[21] ),
    .A2(\sha256cu.m_out_digest.a_in[21] ),
    .B1(_02783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02784_));
 sky130_fd_sc_hd__mux2_2 _08176_ (.A0(\sha256cu.m_out_digest.g_in[21] ),
    .A1(\sha256cu.m_out_digest.f_in[21] ),
    .S(\sha256cu.m_out_digest.e_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02785_));
 sky130_fd_sc_hd__xnor2_1 _08177_ (.A(_02784_),
    .B(_02785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02786_));
 sky130_fd_sc_hd__xor2_1 _08178_ (.A(\sha256cu.iter_processing.w[21] ),
    .B(_02786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02787_));
 sky130_fd_sc_hd__xnor2_1 _08179_ (.A(_02782_),
    .B(_02787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02788_));
 sky130_fd_sc_hd__and2b_1 _08180_ (.A_N(_02750_),
    .B(_02748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02789_));
 sky130_fd_sc_hd__a21oi_1 _08181_ (.A1(_02742_),
    .A2(_02751_),
    .B1(_02789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02790_));
 sky130_fd_sc_hd__xnor2_1 _08182_ (.A(_02788_),
    .B(_02790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02791_));
 sky130_fd_sc_hd__xnor2_1 _08183_ (.A(_02772_),
    .B(_02791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02792_));
 sky130_fd_sc_hd__or2b_1 _08184_ (.A(_02754_),
    .B_N(_02752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02793_));
 sky130_fd_sc_hd__a21bo_1 _08185_ (.A1(_02737_),
    .A2(_02755_),
    .B1_N(_02793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02794_));
 sky130_fd_sc_hd__xnor2_1 _08186_ (.A(_02792_),
    .B(_02794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02795_));
 sky130_fd_sc_hd__or2_1 _08187_ (.A(\sha256cu.K[21] ),
    .B(_02795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02796_));
 sky130_fd_sc_hd__nand2_1 _08188_ (.A(\sha256cu.K[21] ),
    .B(_02795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_1 _08189_ (.A(_02796_),
    .B(_02797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02798_));
 sky130_fd_sc_hd__or2b_1 _08190_ (.A(_02756_),
    .B_N(_02735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02799_));
 sky130_fd_sc_hd__a21boi_2 _08191_ (.A1(\sha256cu.K[20] ),
    .A2(_02757_),
    .B1_N(_02799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02800_));
 sky130_fd_sc_hd__xnor2_1 _08192_ (.A(_02798_),
    .B(_02800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02801_));
 sky130_fd_sc_hd__o22a_1 _08193_ (.A1(_02758_),
    .A2(_02760_),
    .B1(_02761_),
    .B2(_02767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02802_));
 sky130_fd_sc_hd__xor2_1 _08194_ (.A(_02801_),
    .B(_02802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02803_));
 sky130_fd_sc_hd__or2_1 _08195_ (.A(\sha256cu.m_out_digest.a_in[21] ),
    .B(_02440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02804_));
 sky130_fd_sc_hd__o211a_1 _08196_ (.A1(_02332_),
    .A2(_02803_),
    .B1(_02804_),
    .C1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00116_));
 sky130_fd_sc_hd__or2b_1 _08197_ (.A(_02792_),
    .B_N(_02794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02805_));
 sky130_fd_sc_hd__inv_2 _08198_ (.A(\sha256cu.K[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02806_));
 sky130_fd_sc_hd__xnor2_2 _08199_ (.A(_02382_),
    .B(\sha256cu.m_out_digest.a_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02807_));
 sky130_fd_sc_hd__xnor2_1 _08200_ (.A(_02083_),
    .B(_02807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02808_));
 sky130_fd_sc_hd__xnor2_1 _08201_ (.A(\sha256cu.m_out_digest.h_in[22] ),
    .B(_02808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02809_));
 sky130_fd_sc_hd__xnor2_4 _08202_ (.A(\sha256cu.m_out_digest.e_in[15] ),
    .B(\sha256cu.m_out_digest.e_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02810_));
 sky130_fd_sc_hd__xnor2_4 _08203_ (.A(\sha256cu.m_out_digest.e_in[28] ),
    .B(_02810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02811_));
 sky130_fd_sc_hd__xnor2_1 _08204_ (.A(_02809_),
    .B(_02811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02812_));
 sky130_fd_sc_hd__inv_2 _08205_ (.A(_02777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02813_));
 sky130_fd_sc_hd__nand2_1 _08206_ (.A(\sha256cu.m_out_digest.h_in[21] ),
    .B(_02774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02814_));
 sky130_fd_sc_hd__o21a_1 _08207_ (.A1(_02775_),
    .A2(_02813_),
    .B1(_02814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02815_));
 sky130_fd_sc_hd__xnor2_1 _08208_ (.A(_02812_),
    .B(_02815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02816_));
 sky130_fd_sc_hd__a21o_1 _08209_ (.A1(\sha256cu.m_out_digest.b_in[22] ),
    .A2(_02026_),
    .B1(\sha256cu.m_out_digest.c_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02817_));
 sky130_fd_sc_hd__o21ai_1 _08210_ (.A1(\sha256cu.m_out_digest.b_in[22] ),
    .A2(_02026_),
    .B1(_02817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02818_));
 sky130_fd_sc_hd__mux2_2 _08211_ (.A0(\sha256cu.m_out_digest.g_in[22] ),
    .A1(\sha256cu.m_out_digest.f_in[22] ),
    .S(\sha256cu.m_out_digest.e_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02819_));
 sky130_fd_sc_hd__xnor2_1 _08212_ (.A(_02818_),
    .B(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02820_));
 sky130_fd_sc_hd__nor2_1 _08213_ (.A(\sha256cu.iter_processing.w[22] ),
    .B(_02820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02821_));
 sky130_fd_sc_hd__and2_1 _08214_ (.A(\sha256cu.iter_processing.w[22] ),
    .B(_02820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02822_));
 sky130_fd_sc_hd__nor2_1 _08215_ (.A(_02821_),
    .B(_02822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02823_));
 sky130_fd_sc_hd__xnor2_1 _08216_ (.A(_02816_),
    .B(_02823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02824_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_02778_),
    .B(_02781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02825_));
 sky130_fd_sc_hd__a21boi_1 _08218_ (.A1(_02782_),
    .A2(_02787_),
    .B1_N(_02825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02826_));
 sky130_fd_sc_hd__nor2_1 _08219_ (.A(_02824_),
    .B(_02826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02827_));
 sky130_fd_sc_hd__and2_1 _08220_ (.A(_02824_),
    .B(_02826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02828_));
 sky130_fd_sc_hd__or2_1 _08221_ (.A(_02827_),
    .B(_02828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02829_));
 sky130_fd_sc_hd__and2b_1 _08222_ (.A_N(_02784_),
    .B(_02785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02830_));
 sky130_fd_sc_hd__a21oi_1 _08223_ (.A1(\sha256cu.iter_processing.w[21] ),
    .A2(_02786_),
    .B1(_02830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02831_));
 sky130_fd_sc_hd__xnor2_1 _08224_ (.A(_02829_),
    .B(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02832_));
 sky130_fd_sc_hd__or2_1 _08225_ (.A(_02788_),
    .B(_02790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02833_));
 sky130_fd_sc_hd__o21ai_1 _08226_ (.A1(_02772_),
    .A2(_02791_),
    .B1(_02833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02834_));
 sky130_fd_sc_hd__xor2_1 _08227_ (.A(_02832_),
    .B(_02834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02835_));
 sky130_fd_sc_hd__xnor2_1 _08228_ (.A(_02806_),
    .B(_02835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02836_));
 sky130_fd_sc_hd__a21oi_1 _08229_ (.A1(_02805_),
    .A2(_02797_),
    .B1(_02836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02837_));
 sky130_fd_sc_hd__and3_1 _08230_ (.A(_02805_),
    .B(_02797_),
    .C(_02836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02838_));
 sky130_fd_sc_hd__or2_1 _08231_ (.A(_02837_),
    .B(_02838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02839_));
 sky130_fd_sc_hd__or2_1 _08232_ (.A(_02761_),
    .B(_02801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02840_));
 sky130_fd_sc_hd__a211o_1 _08233_ (.A1(_02798_),
    .A2(_02800_),
    .B1(_02758_),
    .C1(_02760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02841_));
 sky130_fd_sc_hd__o21ai_1 _08234_ (.A1(_02798_),
    .A2(_02800_),
    .B1(_02841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02842_));
 sky130_fd_sc_hd__o21ba_1 _08235_ (.A1(_02767_),
    .A2(_02840_),
    .B1_N(_02842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02843_));
 sky130_fd_sc_hd__xnor2_1 _08236_ (.A(_02839_),
    .B(_02843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02844_));
 sky130_fd_sc_hd__nor2_1 _08237_ (.A(_02069_),
    .B(_02844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02845_));
 sky130_fd_sc_hd__a22o_1 _08238_ (.A1(_02026_),
    .A2(_02070_),
    .B1(_02845_),
    .B2(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00117_));
 sky130_fd_sc_hd__and2b_1 _08239_ (.A_N(_02818_),
    .B(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02846_));
 sky130_fd_sc_hd__xnor2_2 _08240_ (.A(_02027_),
    .B(\sha256cu.m_out_digest.a_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02847_));
 sky130_fd_sc_hd__xnor2_1 _08241_ (.A(\sha256cu.m_out_digest.a_in[25] ),
    .B(_02847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02848_));
 sky130_fd_sc_hd__xnor2_1 _08242_ (.A(\sha256cu.m_out_digest.h_in[23] ),
    .B(_02848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02849_));
 sky130_fd_sc_hd__xnor2_4 _08243_ (.A(\sha256cu.m_out_digest.e_in[16] ),
    .B(\sha256cu.m_out_digest.e_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02850_));
 sky130_fd_sc_hd__xnor2_4 _08244_ (.A(\sha256cu.m_out_digest.e_in[29] ),
    .B(_02850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02851_));
 sky130_fd_sc_hd__xnor2_1 _08245_ (.A(_02849_),
    .B(_02851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02852_));
 sky130_fd_sc_hd__or2_1 _08246_ (.A(\sha256cu.m_out_digest.h_in[22] ),
    .B(_02808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02853_));
 sky130_fd_sc_hd__and2_1 _08247_ (.A(\sha256cu.m_out_digest.h_in[22] ),
    .B(_02808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02854_));
 sky130_fd_sc_hd__a21oi_1 _08248_ (.A1(_02853_),
    .A2(_02811_),
    .B1(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02855_));
 sky130_fd_sc_hd__xnor2_1 _08249_ (.A(_02852_),
    .B(_02855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02856_));
 sky130_fd_sc_hd__a21o_1 _08250_ (.A1(\sha256cu.m_out_digest.b_in[23] ),
    .A2(\sha256cu.m_out_digest.a_in[23] ),
    .B1(\sha256cu.m_out_digest.c_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02857_));
 sky130_fd_sc_hd__o21ai_1 _08251_ (.A1(\sha256cu.m_out_digest.b_in[23] ),
    .A2(\sha256cu.m_out_digest.a_in[23] ),
    .B1(_02857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02858_));
 sky130_fd_sc_hd__mux2_2 _08252_ (.A0(\sha256cu.m_out_digest.g_in[23] ),
    .A1(\sha256cu.m_out_digest.f_in[23] ),
    .S(\sha256cu.m_out_digest.e_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02859_));
 sky130_fd_sc_hd__xnor2_1 _08253_ (.A(_02858_),
    .B(_02859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02860_));
 sky130_fd_sc_hd__xor2_1 _08254_ (.A(\sha256cu.iter_processing.w[23] ),
    .B(_02860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02861_));
 sky130_fd_sc_hd__xnor2_1 _08255_ (.A(_02856_),
    .B(_02861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02862_));
 sky130_fd_sc_hd__and2b_1 _08256_ (.A_N(_02815_),
    .B(_02812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02863_));
 sky130_fd_sc_hd__a21oi_1 _08257_ (.A1(_02816_),
    .A2(_02823_),
    .B1(_02863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02864_));
 sky130_fd_sc_hd__xnor2_1 _08258_ (.A(_02862_),
    .B(_02864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02865_));
 sky130_fd_sc_hd__o21ba_1 _08259_ (.A1(_02846_),
    .A2(_02822_),
    .B1_N(_02865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02866_));
 sky130_fd_sc_hd__or3b_1 _08260_ (.A(_02846_),
    .B(_02822_),
    .C_N(_02865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02867_));
 sky130_fd_sc_hd__or2b_1 _08261_ (.A(_02866_),
    .B_N(_02867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02868_));
 sky130_fd_sc_hd__o21bai_1 _08262_ (.A1(_02829_),
    .A2(_02831_),
    .B1_N(_02827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02869_));
 sky130_fd_sc_hd__xnor2_1 _08263_ (.A(_02868_),
    .B(_02869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02870_));
 sky130_fd_sc_hd__xnor2_2 _08264_ (.A(\sha256cu.K[23] ),
    .B(_02870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02871_));
 sky130_fd_sc_hd__or2b_1 _08265_ (.A(_02832_),
    .B_N(_02834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02872_));
 sky130_fd_sc_hd__o21ai_2 _08266_ (.A1(_02806_),
    .A2(_02835_),
    .B1(_02872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02873_));
 sky130_fd_sc_hd__xor2_2 _08267_ (.A(_02871_),
    .B(_02873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02874_));
 sky130_fd_sc_hd__o21bai_1 _08268_ (.A1(_02839_),
    .A2(_02843_),
    .B1_N(_02837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02875_));
 sky130_fd_sc_hd__xnor2_1 _08269_ (.A(_02874_),
    .B(_02875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02876_));
 sky130_fd_sc_hd__or2_1 _08270_ (.A(\sha256cu.m_out_digest.a_in[23] ),
    .B(_02440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02877_));
 sky130_fd_sc_hd__o211a_1 _08271_ (.A1(_02332_),
    .A2(_02876_),
    .B1(_02877_),
    .C1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00118_));
 sky130_fd_sc_hd__or3_1 _08272_ (.A(_02839_),
    .B(_02840_),
    .C(_02874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02878_));
 sky130_fd_sc_hd__a211o_1 _08273_ (.A1(_02623_),
    .A2(_02626_),
    .B1(_02763_),
    .C1(_02878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02879_));
 sky130_fd_sc_hd__or3b_1 _08274_ (.A(_02839_),
    .B(_02874_),
    .C_N(_02842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02880_));
 sky130_fd_sc_hd__or2b_1 _08275_ (.A(_02873_),
    .B_N(_02871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02881_));
 sky130_fd_sc_hd__and2b_1 _08276_ (.A_N(_02871_),
    .B(_02873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02882_));
 sky130_fd_sc_hd__a21oi_1 _08277_ (.A1(_02837_),
    .A2(_02881_),
    .B1(_02882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02883_));
 sky130_fd_sc_hd__o211a_1 _08278_ (.A1(_02766_),
    .A2(_02878_),
    .B1(_02880_),
    .C1(_02883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02884_));
 sky130_fd_sc_hd__and2_1 _08279_ (.A(_02879_),
    .B(_02884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02885_));
 sky130_fd_sc_hd__and2b_1 _08280_ (.A_N(_02868_),
    .B(_02869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02886_));
 sky130_fd_sc_hd__and2_1 _08281_ (.A(\sha256cu.K[23] ),
    .B(_02870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02887_));
 sky130_fd_sc_hd__inv_2 _08282_ (.A(\sha256cu.K[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02888_));
 sky130_fd_sc_hd__or2b_1 _08283_ (.A(_02855_),
    .B_N(_02852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02889_));
 sky130_fd_sc_hd__nand2_1 _08284_ (.A(_02856_),
    .B(_02861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02890_));
 sky130_fd_sc_hd__xnor2_2 _08285_ (.A(\sha256cu.m_out_digest.a_in[14] ),
    .B(\sha256cu.m_out_digest.a_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02891_));
 sky130_fd_sc_hd__xnor2_1 _08286_ (.A(_02161_),
    .B(_02891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02892_));
 sky130_fd_sc_hd__xnor2_1 _08287_ (.A(\sha256cu.m_out_digest.h_in[24] ),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02893_));
 sky130_fd_sc_hd__xnor2_2 _08288_ (.A(\sha256cu.m_out_digest.e_in[17] ),
    .B(\sha256cu.m_out_digest.e_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02894_));
 sky130_fd_sc_hd__xnor2_4 _08289_ (.A(\sha256cu.m_out_digest.e_in[30] ),
    .B(_02894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02895_));
 sky130_fd_sc_hd__xnor2_1 _08290_ (.A(_02893_),
    .B(_02895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02896_));
 sky130_fd_sc_hd__or2_1 _08291_ (.A(\sha256cu.m_out_digest.h_in[23] ),
    .B(_02848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02897_));
 sky130_fd_sc_hd__and2_1 _08292_ (.A(\sha256cu.m_out_digest.h_in[23] ),
    .B(_02848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02898_));
 sky130_fd_sc_hd__a21oi_1 _08293_ (.A1(_02897_),
    .A2(_02851_),
    .B1(_02898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02899_));
 sky130_fd_sc_hd__xnor2_1 _08294_ (.A(_02896_),
    .B(_02899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02900_));
 sky130_fd_sc_hd__a21o_1 _08295_ (.A1(\sha256cu.m_out_digest.b_in[24] ),
    .A2(_02083_),
    .B1(\sha256cu.m_out_digest.c_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02901_));
 sky130_fd_sc_hd__o21ai_1 _08296_ (.A1(\sha256cu.m_out_digest.b_in[24] ),
    .A2(_02083_),
    .B1(_02901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02902_));
 sky130_fd_sc_hd__mux2_2 _08297_ (.A0(\sha256cu.m_out_digest.g_in[24] ),
    .A1(\sha256cu.m_out_digest.f_in[24] ),
    .S(\sha256cu.m_out_digest.e_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02903_));
 sky130_fd_sc_hd__xnor2_1 _08298_ (.A(_02902_),
    .B(_02903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02904_));
 sky130_fd_sc_hd__xor2_1 _08299_ (.A(\sha256cu.iter_processing.w[24] ),
    .B(_02904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02905_));
 sky130_fd_sc_hd__xnor2_1 _08300_ (.A(_02900_),
    .B(_02905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02906_));
 sky130_fd_sc_hd__a21oi_1 _08301_ (.A1(_02889_),
    .A2(_02890_),
    .B1(_02906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02907_));
 sky130_fd_sc_hd__and3_1 _08302_ (.A(_02889_),
    .B(_02890_),
    .C(_02906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02908_));
 sky130_fd_sc_hd__or2_1 _08303_ (.A(_02907_),
    .B(_02908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02909_));
 sky130_fd_sc_hd__and2b_1 _08304_ (.A_N(_02858_),
    .B(_02859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02910_));
 sky130_fd_sc_hd__a21oi_1 _08305_ (.A1(\sha256cu.iter_processing.w[23] ),
    .A2(_02860_),
    .B1(_02910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02911_));
 sky130_fd_sc_hd__xnor2_1 _08306_ (.A(_02909_),
    .B(_02911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02912_));
 sky130_fd_sc_hd__o21ba_1 _08307_ (.A1(_02862_),
    .A2(_02864_),
    .B1_N(_02866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02913_));
 sky130_fd_sc_hd__or2_1 _08308_ (.A(_02912_),
    .B(_02913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02914_));
 sky130_fd_sc_hd__nand2_1 _08309_ (.A(_02912_),
    .B(_02913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02915_));
 sky130_fd_sc_hd__nand2_1 _08310_ (.A(_02914_),
    .B(_02915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02916_));
 sky130_fd_sc_hd__xnor2_1 _08311_ (.A(_02888_),
    .B(_02916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02917_));
 sky130_fd_sc_hd__o21ba_1 _08312_ (.A1(_02886_),
    .A2(_02887_),
    .B1_N(_02917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02918_));
 sky130_fd_sc_hd__or3b_1 _08313_ (.A(_02886_),
    .B(_02887_),
    .C_N(_02917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02919_));
 sky130_fd_sc_hd__or2b_2 _08314_ (.A(_02918_),
    .B_N(_02919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02920_));
 sky130_fd_sc_hd__or2_1 _08315_ (.A(_02885_),
    .B(_02920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02921_));
 sky130_fd_sc_hd__nand2_1 _08316_ (.A(_02885_),
    .B(_02920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02922_));
 sky130_fd_sc_hd__a32o_1 _08317_ (.A1(_02113_),
    .A2(_02921_),
    .A3(_02922_),
    .B1(_02332_),
    .B2(_02083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00119_));
 sky130_fd_sc_hd__clkbuf_4 _08318_ (.A(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02923_));
 sky130_fd_sc_hd__inv_2 _08319_ (.A(\sha256cu.K[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02924_));
 sky130_fd_sc_hd__or2b_1 _08320_ (.A(_02899_),
    .B_N(_02896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02925_));
 sky130_fd_sc_hd__nand2_1 _08321_ (.A(_02900_),
    .B(_02905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02926_));
 sky130_fd_sc_hd__xnor2_2 _08322_ (.A(_02084_),
    .B(\sha256cu.m_out_digest.a_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02927_));
 sky130_fd_sc_hd__xnor2_1 _08323_ (.A(\sha256cu.m_out_digest.a_in[27] ),
    .B(_02927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02928_));
 sky130_fd_sc_hd__xnor2_1 _08324_ (.A(\sha256cu.m_out_digest.h_in[25] ),
    .B(_02928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02929_));
 sky130_fd_sc_hd__xnor2_4 _08325_ (.A(\sha256cu.m_out_digest.e_in[18] ),
    .B(\sha256cu.m_out_digest.e_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02930_));
 sky130_fd_sc_hd__xnor2_4 _08326_ (.A(\sha256cu.m_out_digest.e_in[31] ),
    .B(_02930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02931_));
 sky130_fd_sc_hd__xnor2_1 _08327_ (.A(_02929_),
    .B(_02931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02932_));
 sky130_fd_sc_hd__or2_1 _08328_ (.A(\sha256cu.m_out_digest.h_in[24] ),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02933_));
 sky130_fd_sc_hd__and2_1 _08329_ (.A(\sha256cu.m_out_digest.h_in[24] ),
    .B(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02934_));
 sky130_fd_sc_hd__a21o_1 _08330_ (.A1(_02933_),
    .A2(_02895_),
    .B1(_02934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02935_));
 sky130_fd_sc_hd__xor2_1 _08331_ (.A(_02932_),
    .B(_02935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02936_));
 sky130_fd_sc_hd__a21o_1 _08332_ (.A1(\sha256cu.m_out_digest.b_in[25] ),
    .A2(\sha256cu.m_out_digest.a_in[25] ),
    .B1(\sha256cu.m_out_digest.c_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02937_));
 sky130_fd_sc_hd__o21ai_1 _08333_ (.A1(\sha256cu.m_out_digest.b_in[25] ),
    .A2(\sha256cu.m_out_digest.a_in[25] ),
    .B1(_02937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02938_));
 sky130_fd_sc_hd__mux2_1 _08334_ (.A0(\sha256cu.m_out_digest.g_in[25] ),
    .A1(\sha256cu.m_out_digest.f_in[25] ),
    .S(\sha256cu.m_out_digest.e_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02939_));
 sky130_fd_sc_hd__xnor2_1 _08335_ (.A(_02938_),
    .B(_02939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02940_));
 sky130_fd_sc_hd__xor2_1 _08336_ (.A(\sha256cu.iter_processing.w[25] ),
    .B(_02940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02941_));
 sky130_fd_sc_hd__xnor2_1 _08337_ (.A(_02936_),
    .B(_02941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02942_));
 sky130_fd_sc_hd__a21oi_1 _08338_ (.A1(_02925_),
    .A2(_02926_),
    .B1(_02942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02943_));
 sky130_fd_sc_hd__and3_1 _08339_ (.A(_02925_),
    .B(_02926_),
    .C(_02942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02944_));
 sky130_fd_sc_hd__or2_1 _08340_ (.A(_02943_),
    .B(_02944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02945_));
 sky130_fd_sc_hd__and2b_1 _08341_ (.A_N(_02902_),
    .B(_02903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02946_));
 sky130_fd_sc_hd__a21oi_1 _08342_ (.A1(\sha256cu.iter_processing.w[24] ),
    .A2(_02904_),
    .B1(_02946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02947_));
 sky130_fd_sc_hd__xnor2_1 _08343_ (.A(_02945_),
    .B(_02947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02948_));
 sky130_fd_sc_hd__o21ba_1 _08344_ (.A1(_02909_),
    .A2(_02911_),
    .B1_N(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02949_));
 sky130_fd_sc_hd__xnor2_1 _08345_ (.A(_02948_),
    .B(_02949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02950_));
 sky130_fd_sc_hd__and2_1 _08346_ (.A(_02924_),
    .B(_02950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02951_));
 sky130_fd_sc_hd__nor2_1 _08347_ (.A(_02924_),
    .B(_02950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02952_));
 sky130_fd_sc_hd__or2_1 _08348_ (.A(_02951_),
    .B(_02952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02953_));
 sky130_fd_sc_hd__o21a_1 _08349_ (.A1(_02888_),
    .A2(_02916_),
    .B1(_02914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02954_));
 sky130_fd_sc_hd__xnor2_1 _08350_ (.A(_02953_),
    .B(_02954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02955_));
 sky130_fd_sc_hd__o21ba_1 _08351_ (.A1(_02885_),
    .A2(_02920_),
    .B1_N(_02918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02956_));
 sky130_fd_sc_hd__xnor2_1 _08352_ (.A(_02955_),
    .B(_02956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02957_));
 sky130_fd_sc_hd__o2bb2a_1 _08353_ (.A1_N(\sha256cu.m_out_digest.a_in[25] ),
    .A2_N(_02629_),
    .B1(_02923_),
    .B2(_02957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02958_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_02000_),
    .B(_02958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00120_));
 sky130_fd_sc_hd__nor2_1 _08355_ (.A(_02945_),
    .B(_02947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02959_));
 sky130_fd_sc_hd__xnor2_1 _08356_ (.A(_02128_),
    .B(\sha256cu.m_out_digest.a_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02960_));
 sky130_fd_sc_hd__xnor2_1 _08357_ (.A(_02232_),
    .B(_02960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02961_));
 sky130_fd_sc_hd__xnor2_1 _08358_ (.A(\sha256cu.m_out_digest.h_in[26] ),
    .B(_02961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02962_));
 sky130_fd_sc_hd__xnor2_2 _08359_ (.A(\sha256cu.m_out_digest.e_in[5] ),
    .B(\sha256cu.m_out_digest.e_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02963_));
 sky130_fd_sc_hd__xnor2_4 _08360_ (.A(\sha256cu.m_out_digest.e_in[19] ),
    .B(_02963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02964_));
 sky130_fd_sc_hd__xnor2_1 _08361_ (.A(_02962_),
    .B(_02964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02965_));
 sky130_fd_sc_hd__and2b_1 _08362_ (.A_N(_02929_),
    .B(_02931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02966_));
 sky130_fd_sc_hd__a21oi_1 _08363_ (.A1(\sha256cu.m_out_digest.h_in[25] ),
    .A2(_02928_),
    .B1(_02966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02967_));
 sky130_fd_sc_hd__xnor2_1 _08364_ (.A(_02965_),
    .B(_02967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02968_));
 sky130_fd_sc_hd__a21o_1 _08365_ (.A1(\sha256cu.m_out_digest.b_in[26] ),
    .A2(_02161_),
    .B1(\sha256cu.m_out_digest.c_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02969_));
 sky130_fd_sc_hd__o21ai_1 _08366_ (.A1(\sha256cu.m_out_digest.b_in[26] ),
    .A2(_02161_),
    .B1(_02969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02970_));
 sky130_fd_sc_hd__mux2_2 _08367_ (.A0(\sha256cu.m_out_digest.g_in[26] ),
    .A1(\sha256cu.m_out_digest.f_in[26] ),
    .S(\sha256cu.m_out_digest.e_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02971_));
 sky130_fd_sc_hd__xnor2_1 _08368_ (.A(_02970_),
    .B(_02971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02972_));
 sky130_fd_sc_hd__xor2_1 _08369_ (.A(\sha256cu.iter_processing.w[26] ),
    .B(_02972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02973_));
 sky130_fd_sc_hd__xnor2_1 _08370_ (.A(_02968_),
    .B(_02973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_1 _08371_ (.A(_02932_),
    .B(_02935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02975_));
 sky130_fd_sc_hd__a21bo_1 _08372_ (.A1(_02936_),
    .A2(_02941_),
    .B1_N(_02975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02976_));
 sky130_fd_sc_hd__xor2_1 _08373_ (.A(_02974_),
    .B(_02976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02977_));
 sky130_fd_sc_hd__and2b_1 _08374_ (.A_N(_02938_),
    .B(_02939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02978_));
 sky130_fd_sc_hd__a21oi_1 _08375_ (.A1(\sha256cu.iter_processing.w[25] ),
    .A2(_02940_),
    .B1(_02978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02979_));
 sky130_fd_sc_hd__xnor2_1 _08376_ (.A(_02977_),
    .B(_02979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02980_));
 sky130_fd_sc_hd__o21ba_1 _08377_ (.A1(_02943_),
    .A2(_02959_),
    .B1_N(_02980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02981_));
 sky130_fd_sc_hd__or3b_1 _08378_ (.A(_02943_),
    .B(_02959_),
    .C_N(_02980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02982_));
 sky130_fd_sc_hd__or2b_1 _08379_ (.A(_02981_),
    .B_N(_02982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02983_));
 sky130_fd_sc_hd__and2b_1 _08380_ (.A_N(\sha256cu.K[26] ),
    .B(_02983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02984_));
 sky130_fd_sc_hd__and3b_1 _08381_ (.A_N(_02981_),
    .B(_02982_),
    .C(\sha256cu.K[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02985_));
 sky130_fd_sc_hd__or2_1 _08382_ (.A(_02984_),
    .B(_02985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02986_));
 sky130_fd_sc_hd__o21ba_1 _08383_ (.A1(_02948_),
    .A2(_02949_),
    .B1_N(_02952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02987_));
 sky130_fd_sc_hd__xnor2_2 _08384_ (.A(_02986_),
    .B(_02987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02988_));
 sky130_fd_sc_hd__or2_1 _08385_ (.A(_02920_),
    .B(_02955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02989_));
 sky130_fd_sc_hd__nor2_1 _08386_ (.A(_02953_),
    .B(_02954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02990_));
 sky130_fd_sc_hd__nand2_1 _08387_ (.A(_02953_),
    .B(_02954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02991_));
 sky130_fd_sc_hd__o21a_1 _08388_ (.A1(_02918_),
    .A2(_02990_),
    .B1(_02991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02992_));
 sky130_fd_sc_hd__o21ba_1 _08389_ (.A1(_02885_),
    .A2(_02989_),
    .B1_N(_02992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02993_));
 sky130_fd_sc_hd__nor2_1 _08390_ (.A(_02988_),
    .B(_02993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02994_));
 sky130_fd_sc_hd__a21o_1 _08391_ (.A1(_02988_),
    .A2(_02993_),
    .B1(_02478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02995_));
 sky130_fd_sc_hd__a2bb2o_1 _08392_ (.A1_N(_02994_),
    .A2_N(_02995_),
    .B1(_02161_),
    .B2(_02070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00121_));
 sky130_fd_sc_hd__inv_2 _08393_ (.A(\sha256cu.K[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02996_));
 sky130_fd_sc_hd__xnor2_1 _08394_ (.A(_02162_),
    .B(\sha256cu.m_out_digest.a_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02997_));
 sky130_fd_sc_hd__xnor2_1 _08395_ (.A(_02272_),
    .B(_02997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02998_));
 sky130_fd_sc_hd__xnor2_1 _08396_ (.A(\sha256cu.m_out_digest.h_in[27] ),
    .B(_02998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02999_));
 sky130_fd_sc_hd__xnor2_4 _08397_ (.A(\sha256cu.m_out_digest.e_in[6] ),
    .B(\sha256cu.m_out_digest.e_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03000_));
 sky130_fd_sc_hd__xnor2_4 _08398_ (.A(\sha256cu.m_out_digest.e_in[20] ),
    .B(_03000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03001_));
 sky130_fd_sc_hd__xnor2_1 _08399_ (.A(_02999_),
    .B(_03001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03002_));
 sky130_fd_sc_hd__or2b_1 _08400_ (.A(_02962_),
    .B_N(_02964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03003_));
 sky130_fd_sc_hd__a21bo_1 _08401_ (.A1(\sha256cu.m_out_digest.h_in[26] ),
    .A2(_02961_),
    .B1_N(_03003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03004_));
 sky130_fd_sc_hd__xor2_1 _08402_ (.A(_03002_),
    .B(_03004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03005_));
 sky130_fd_sc_hd__a21o_1 _08403_ (.A1(\sha256cu.m_out_digest.b_in[27] ),
    .A2(\sha256cu.m_out_digest.a_in[27] ),
    .B1(\sha256cu.m_out_digest.c_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03006_));
 sky130_fd_sc_hd__o21ai_1 _08404_ (.A1(\sha256cu.m_out_digest.b_in[27] ),
    .A2(\sha256cu.m_out_digest.a_in[27] ),
    .B1(_03006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03007_));
 sky130_fd_sc_hd__mux2_1 _08405_ (.A0(\sha256cu.m_out_digest.g_in[27] ),
    .A1(\sha256cu.m_out_digest.f_in[27] ),
    .S(\sha256cu.m_out_digest.e_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03008_));
 sky130_fd_sc_hd__xnor2_1 _08406_ (.A(_03007_),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03009_));
 sky130_fd_sc_hd__xor2_1 _08407_ (.A(\sha256cu.iter_processing.w[27] ),
    .B(_03009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03010_));
 sky130_fd_sc_hd__nand2_1 _08408_ (.A(_03005_),
    .B(_03010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03011_));
 sky130_fd_sc_hd__or2_1 _08409_ (.A(_03005_),
    .B(_03010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03012_));
 sky130_fd_sc_hd__nand2_1 _08410_ (.A(_03011_),
    .B(_03012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03013_));
 sky130_fd_sc_hd__or2b_1 _08411_ (.A(_02967_),
    .B_N(_02965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03014_));
 sky130_fd_sc_hd__a21bo_1 _08412_ (.A1(_02968_),
    .A2(_02973_),
    .B1_N(_03014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03015_));
 sky130_fd_sc_hd__xor2_1 _08413_ (.A(_03013_),
    .B(_03015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03016_));
 sky130_fd_sc_hd__and2b_1 _08414_ (.A_N(_02970_),
    .B(_02971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03017_));
 sky130_fd_sc_hd__a21oi_1 _08415_ (.A1(\sha256cu.iter_processing.w[26] ),
    .A2(_02972_),
    .B1(_03017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03018_));
 sky130_fd_sc_hd__xnor2_1 _08416_ (.A(_03016_),
    .B(_03018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03019_));
 sky130_fd_sc_hd__and2b_1 _08417_ (.A_N(_02974_),
    .B(_02976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03020_));
 sky130_fd_sc_hd__o21ba_1 _08418_ (.A1(_02977_),
    .A2(_02979_),
    .B1_N(_03020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03021_));
 sky130_fd_sc_hd__xnor2_1 _08419_ (.A(_03019_),
    .B(_03021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03022_));
 sky130_fd_sc_hd__xnor2_1 _08420_ (.A(_02996_),
    .B(_03022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03023_));
 sky130_fd_sc_hd__o21ba_1 _08421_ (.A1(_02981_),
    .A2(_02985_),
    .B1_N(_03023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03024_));
 sky130_fd_sc_hd__or3b_1 _08422_ (.A(_02981_),
    .B(_02985_),
    .C_N(_03023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03025_));
 sky130_fd_sc_hd__nand2b_1 _08423_ (.A_N(_03024_),
    .B(_03025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03026_));
 sky130_fd_sc_hd__nor2_1 _08424_ (.A(_02986_),
    .B(_02987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03027_));
 sky130_fd_sc_hd__o21ba_1 _08425_ (.A1(_02988_),
    .A2(_02993_),
    .B1_N(_03027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03028_));
 sky130_fd_sc_hd__xor2_1 _08426_ (.A(_03026_),
    .B(_03028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03029_));
 sky130_fd_sc_hd__and2_1 _08427_ (.A(\sha256cu.m_out_digest.a_in[27] ),
    .B(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03030_));
 sky130_fd_sc_hd__a211o_1 _08428_ (.A1(_02369_),
    .A2(_03029_),
    .B1(_03030_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00122_));
 sky130_fd_sc_hd__clkbuf_8 _08429_ (.A(_02069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03031_));
 sky130_fd_sc_hd__nor2_1 _08430_ (.A(_02988_),
    .B(_03026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03032_));
 sky130_fd_sc_hd__a221oi_2 _08431_ (.A1(_03027_),
    .A2(_03025_),
    .B1(_03032_),
    .B2(_02992_),
    .C1(_03024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03033_));
 sky130_fd_sc_hd__a2111o_1 _08432_ (.A1(_02879_),
    .A2(_02884_),
    .B1(_02988_),
    .C1(_02989_),
    .D1(_03026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03034_));
 sky130_fd_sc_hd__nor2_1 _08433_ (.A(_03019_),
    .B(_03021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03035_));
 sky130_fd_sc_hd__nor2_1 _08434_ (.A(_02996_),
    .B(_03022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03036_));
 sky130_fd_sc_hd__inv_2 _08435_ (.A(\sha256cu.K[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03037_));
 sky130_fd_sc_hd__and3_1 _08436_ (.A(_03011_),
    .B(_03012_),
    .C(_03015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03038_));
 sky130_fd_sc_hd__nor2_1 _08437_ (.A(_03016_),
    .B(_03018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03039_));
 sky130_fd_sc_hd__nand2_1 _08438_ (.A(_03002_),
    .B(_03004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03040_));
 sky130_fd_sc_hd__xnor2_1 _08439_ (.A(_02198_),
    .B(\sha256cu.m_out_digest.a_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03041_));
 sky130_fd_sc_hd__xnor2_2 _08440_ (.A(_02304_),
    .B(_03041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03042_));
 sky130_fd_sc_hd__xnor2_1 _08441_ (.A(\sha256cu.m_out_digest.h_in[28] ),
    .B(_03042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03043_));
 sky130_fd_sc_hd__xnor2_4 _08442_ (.A(\sha256cu.m_out_digest.e_in[7] ),
    .B(\sha256cu.m_out_digest.e_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03044_));
 sky130_fd_sc_hd__xnor2_4 _08443_ (.A(\sha256cu.m_out_digest.e_in[21] ),
    .B(_03044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03045_));
 sky130_fd_sc_hd__xnor2_1 _08444_ (.A(_03043_),
    .B(_03045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03046_));
 sky130_fd_sc_hd__or2b_1 _08445_ (.A(_02999_),
    .B_N(_03001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03047_));
 sky130_fd_sc_hd__a21bo_1 _08446_ (.A1(\sha256cu.m_out_digest.h_in[27] ),
    .A2(_02998_),
    .B1_N(_03047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03048_));
 sky130_fd_sc_hd__xor2_1 _08447_ (.A(_03046_),
    .B(_03048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03049_));
 sky130_fd_sc_hd__a21o_1 _08448_ (.A1(\sha256cu.m_out_digest.b_in[28] ),
    .A2(_02232_),
    .B1(\sha256cu.m_out_digest.c_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03050_));
 sky130_fd_sc_hd__o21ai_1 _08449_ (.A1(\sha256cu.m_out_digest.b_in[28] ),
    .A2(_02232_),
    .B1(_03050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03051_));
 sky130_fd_sc_hd__mux2_2 _08450_ (.A0(\sha256cu.m_out_digest.g_in[28] ),
    .A1(\sha256cu.m_out_digest.f_in[28] ),
    .S(\sha256cu.m_out_digest.e_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03052_));
 sky130_fd_sc_hd__xnor2_1 _08451_ (.A(_03051_),
    .B(_03052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03053_));
 sky130_fd_sc_hd__xor2_1 _08452_ (.A(\sha256cu.iter_processing.w[28] ),
    .B(_03053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03054_));
 sky130_fd_sc_hd__nand2_1 _08453_ (.A(_03049_),
    .B(_03054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03055_));
 sky130_fd_sc_hd__or2_1 _08454_ (.A(_03049_),
    .B(_03054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03056_));
 sky130_fd_sc_hd__nand2_1 _08455_ (.A(_03055_),
    .B(_03056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03057_));
 sky130_fd_sc_hd__a21oi_1 _08456_ (.A1(_03040_),
    .A2(_03011_),
    .B1(_03057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03058_));
 sky130_fd_sc_hd__and3_1 _08457_ (.A(_03040_),
    .B(_03011_),
    .C(_03057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03059_));
 sky130_fd_sc_hd__or2_1 _08458_ (.A(_03058_),
    .B(_03059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03060_));
 sky130_fd_sc_hd__and2b_1 _08459_ (.A_N(_03007_),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03061_));
 sky130_fd_sc_hd__a21oi_1 _08460_ (.A1(\sha256cu.iter_processing.w[27] ),
    .A2(_03009_),
    .B1(_03061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03062_));
 sky130_fd_sc_hd__xnor2_1 _08461_ (.A(_03060_),
    .B(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03063_));
 sky130_fd_sc_hd__o21bai_1 _08462_ (.A1(_03038_),
    .A2(_03039_),
    .B1_N(_03063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03064_));
 sky130_fd_sc_hd__or3b_1 _08463_ (.A(_03038_),
    .B(_03039_),
    .C_N(_03063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03065_));
 sky130_fd_sc_hd__nand2_1 _08464_ (.A(_03064_),
    .B(_03065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03066_));
 sky130_fd_sc_hd__xnor2_1 _08465_ (.A(_03037_),
    .B(_03066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03067_));
 sky130_fd_sc_hd__o21bai_2 _08466_ (.A1(_03035_),
    .A2(_03036_),
    .B1_N(_03067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03068_));
 sky130_fd_sc_hd__or3b_1 _08467_ (.A(_03035_),
    .B(_03036_),
    .C_N(_03067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03069_));
 sky130_fd_sc_hd__nand2_1 _08468_ (.A(_03068_),
    .B(_03069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03070_));
 sky130_fd_sc_hd__a21o_1 _08469_ (.A1(_03033_),
    .A2(_03034_),
    .B1(_03070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03071_));
 sky130_fd_sc_hd__and3_1 _08470_ (.A(_03070_),
    .B(_03033_),
    .C(_03034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03072_));
 sky130_fd_sc_hd__nor2_1 _08471_ (.A(_02478_),
    .B(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03073_));
 sky130_fd_sc_hd__a22o_1 _08472_ (.A1(_02232_),
    .A2(_03031_),
    .B1(_03071_),
    .B2(_03073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00123_));
 sky130_fd_sc_hd__or2_1 _08473_ (.A(_03037_),
    .B(_03066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03074_));
 sky130_fd_sc_hd__clkinv_2 _08474_ (.A(\sha256cu.K[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03075_));
 sky130_fd_sc_hd__nor2_1 _08475_ (.A(_03060_),
    .B(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03076_));
 sky130_fd_sc_hd__nand2_1 _08476_ (.A(_03046_),
    .B(_03048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03077_));
 sky130_fd_sc_hd__xnor2_1 _08477_ (.A(_02233_),
    .B(\sha256cu.m_out_digest.a_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03078_));
 sky130_fd_sc_hd__xnor2_2 _08478_ (.A(\sha256cu.m_out_digest.a_in[31] ),
    .B(_03078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03079_));
 sky130_fd_sc_hd__xnor2_1 _08479_ (.A(\sha256cu.m_out_digest.h_in[29] ),
    .B(_03079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03080_));
 sky130_fd_sc_hd__xnor2_4 _08480_ (.A(\sha256cu.m_out_digest.e_in[8] ),
    .B(\sha256cu.m_out_digest.e_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03081_));
 sky130_fd_sc_hd__xnor2_4 _08481_ (.A(\sha256cu.m_out_digest.e_in[22] ),
    .B(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03082_));
 sky130_fd_sc_hd__xnor2_1 _08482_ (.A(_03080_),
    .B(_03082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03083_));
 sky130_fd_sc_hd__or2b_1 _08483_ (.A(_03043_),
    .B_N(_03045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03084_));
 sky130_fd_sc_hd__a21bo_1 _08484_ (.A1(\sha256cu.m_out_digest.h_in[28] ),
    .A2(_03042_),
    .B1_N(_03084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03085_));
 sky130_fd_sc_hd__xor2_1 _08485_ (.A(_03083_),
    .B(_03085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03086_));
 sky130_fd_sc_hd__a21o_1 _08486_ (.A1(\sha256cu.m_out_digest.b_in[29] ),
    .A2(_02272_),
    .B1(\sha256cu.m_out_digest.c_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03087_));
 sky130_fd_sc_hd__o21ai_2 _08487_ (.A1(\sha256cu.m_out_digest.b_in[29] ),
    .A2(_02272_),
    .B1(_03087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03088_));
 sky130_fd_sc_hd__mux2_2 _08488_ (.A0(\sha256cu.m_out_digest.g_in[29] ),
    .A1(\sha256cu.m_out_digest.f_in[29] ),
    .S(\sha256cu.m_out_digest.e_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03089_));
 sky130_fd_sc_hd__xnor2_1 _08489_ (.A(_03088_),
    .B(_03089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03090_));
 sky130_fd_sc_hd__xor2_1 _08490_ (.A(\sha256cu.iter_processing.w[29] ),
    .B(_03090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03091_));
 sky130_fd_sc_hd__nand2_1 _08491_ (.A(_03086_),
    .B(_03091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03092_));
 sky130_fd_sc_hd__or2_1 _08492_ (.A(_03086_),
    .B(_03091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03093_));
 sky130_fd_sc_hd__nand2_1 _08493_ (.A(_03092_),
    .B(_03093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03094_));
 sky130_fd_sc_hd__a21oi_1 _08494_ (.A1(_03077_),
    .A2(_03055_),
    .B1(_03094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03095_));
 sky130_fd_sc_hd__and3_1 _08495_ (.A(_03077_),
    .B(_03055_),
    .C(_03094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03096_));
 sky130_fd_sc_hd__or2_1 _08496_ (.A(_03095_),
    .B(_03096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03097_));
 sky130_fd_sc_hd__and2b_1 _08497_ (.A_N(_03051_),
    .B(_03052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03098_));
 sky130_fd_sc_hd__a21oi_1 _08498_ (.A1(\sha256cu.iter_processing.w[28] ),
    .A2(_03053_),
    .B1(_03098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03099_));
 sky130_fd_sc_hd__xnor2_1 _08499_ (.A(_03097_),
    .B(_03099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03100_));
 sky130_fd_sc_hd__o21ba_1 _08500_ (.A1(_03058_),
    .A2(_03076_),
    .B1_N(_03100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03101_));
 sky130_fd_sc_hd__or3b_1 _08501_ (.A(_03058_),
    .B(_03076_),
    .C_N(_03100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03102_));
 sky130_fd_sc_hd__or2b_1 _08502_ (.A(_03101_),
    .B_N(_03102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03103_));
 sky130_fd_sc_hd__xnor2_1 _08503_ (.A(_03075_),
    .B(_03103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03104_));
 sky130_fd_sc_hd__a21o_1 _08504_ (.A1(_03064_),
    .A2(_03074_),
    .B1(_03104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03105_));
 sky130_fd_sc_hd__and3_1 _08505_ (.A(_03064_),
    .B(_03074_),
    .C(_03104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03106_));
 sky130_fd_sc_hd__inv_2 _08506_ (.A(_03106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03107_));
 sky130_fd_sc_hd__nand2_1 _08507_ (.A(_03105_),
    .B(_03107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03108_));
 sky130_fd_sc_hd__nand3_1 _08508_ (.A(_03068_),
    .B(_03071_),
    .C(_03108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03109_));
 sky130_fd_sc_hd__a21oi_1 _08509_ (.A1(_03068_),
    .A2(_03071_),
    .B1(_03108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03110_));
 sky130_fd_sc_hd__nor2_1 _08510_ (.A(_02069_),
    .B(_03110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03111_));
 sky130_fd_sc_hd__a221o_1 _08511_ (.A1(_02272_),
    .A2(_02220_),
    .B1(_03109_),
    .B2(_03111_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00124_));
 sky130_fd_sc_hd__nor2_1 _08512_ (.A(_03075_),
    .B(_03103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03112_));
 sky130_fd_sc_hd__nor2_1 _08513_ (.A(_03097_),
    .B(_03099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _08514_ (.A(_03083_),
    .B(_03085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03114_));
 sky130_fd_sc_hd__xnor2_1 _08515_ (.A(\sha256cu.m_out_digest.a_in[11] ),
    .B(\sha256cu.m_out_digest.a_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03115_));
 sky130_fd_sc_hd__xnor2_2 _08516_ (.A(_02273_),
    .B(_03115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03116_));
 sky130_fd_sc_hd__xnor2_1 _08517_ (.A(\sha256cu.m_out_digest.h_in[30] ),
    .B(_03116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03117_));
 sky130_fd_sc_hd__xnor2_4 _08518_ (.A(\sha256cu.m_out_digest.e_in[9] ),
    .B(\sha256cu.m_out_digest.e_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03118_));
 sky130_fd_sc_hd__xnor2_4 _08519_ (.A(\sha256cu.m_out_digest.e_in[23] ),
    .B(_03118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03119_));
 sky130_fd_sc_hd__xnor2_1 _08520_ (.A(_03117_),
    .B(_03119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03120_));
 sky130_fd_sc_hd__or2b_1 _08521_ (.A(_03080_),
    .B_N(_03082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03121_));
 sky130_fd_sc_hd__a21bo_1 _08522_ (.A1(\sha256cu.m_out_digest.h_in[29] ),
    .A2(_03079_),
    .B1_N(_03121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03122_));
 sky130_fd_sc_hd__xor2_1 _08523_ (.A(_03120_),
    .B(_03122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03123_));
 sky130_fd_sc_hd__a21o_1 _08524_ (.A1(\sha256cu.m_out_digest.b_in[30] ),
    .A2(_02304_),
    .B1(\sha256cu.m_out_digest.c_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03124_));
 sky130_fd_sc_hd__o21ai_1 _08525_ (.A1(\sha256cu.m_out_digest.b_in[30] ),
    .A2(_02304_),
    .B1(_03124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03125_));
 sky130_fd_sc_hd__mux2_2 _08526_ (.A0(\sha256cu.m_out_digest.g_in[30] ),
    .A1(\sha256cu.m_out_digest.f_in[30] ),
    .S(\sha256cu.m_out_digest.e_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03126_));
 sky130_fd_sc_hd__xnor2_1 _08527_ (.A(_03125_),
    .B(_03126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03127_));
 sky130_fd_sc_hd__xor2_1 _08528_ (.A(\sha256cu.iter_processing.w[30] ),
    .B(_03127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03128_));
 sky130_fd_sc_hd__and2_1 _08529_ (.A(_03123_),
    .B(_03128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03129_));
 sky130_fd_sc_hd__nor2_1 _08530_ (.A(_03123_),
    .B(_03128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03130_));
 sky130_fd_sc_hd__or2_1 _08531_ (.A(_03129_),
    .B(_03130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03131_));
 sky130_fd_sc_hd__a21o_1 _08532_ (.A1(_03114_),
    .A2(_03092_),
    .B1(_03131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03132_));
 sky130_fd_sc_hd__nand3_1 _08533_ (.A(_03114_),
    .B(_03092_),
    .C(_03131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03133_));
 sky130_fd_sc_hd__nand2_1 _08534_ (.A(_03132_),
    .B(_03133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03134_));
 sky130_fd_sc_hd__and2b_1 _08535_ (.A_N(_03088_),
    .B(_03089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03135_));
 sky130_fd_sc_hd__a21oi_1 _08536_ (.A1(\sha256cu.iter_processing.w[29] ),
    .A2(_03090_),
    .B1(_03135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03136_));
 sky130_fd_sc_hd__xnor2_1 _08537_ (.A(_03134_),
    .B(_03136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03137_));
 sky130_fd_sc_hd__o21ba_1 _08538_ (.A1(_03095_),
    .A2(_03113_),
    .B1_N(_03137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03138_));
 sky130_fd_sc_hd__or3b_1 _08539_ (.A(_03095_),
    .B(_03113_),
    .C_N(_03137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03139_));
 sky130_fd_sc_hd__or2b_1 _08540_ (.A(_03138_),
    .B_N(_03139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03140_));
 sky130_fd_sc_hd__xor2_1 _08541_ (.A(\sha256cu.K[30] ),
    .B(_03140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03141_));
 sky130_fd_sc_hd__o21bai_1 _08542_ (.A1(_03101_),
    .A2(_03112_),
    .B1_N(_03141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03142_));
 sky130_fd_sc_hd__or3b_1 _08543_ (.A(_03101_),
    .B(_03112_),
    .C_N(_03141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03143_));
 sky130_fd_sc_hd__nand2_1 _08544_ (.A(_03142_),
    .B(_03143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03144_));
 sky130_fd_sc_hd__a311o_1 _08545_ (.A1(_03068_),
    .A2(_03071_),
    .A3(_03105_),
    .B1(_03106_),
    .C1(_03144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03145_));
 sky130_fd_sc_hd__a31o_1 _08546_ (.A1(_03068_),
    .A2(_03071_),
    .A3(_03105_),
    .B1(_03106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03146_));
 sky130_fd_sc_hd__a21oi_1 _08547_ (.A1(_03144_),
    .A2(_03146_),
    .B1(_02069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03147_));
 sky130_fd_sc_hd__a221o_1 _08548_ (.A1(_02304_),
    .A2(_02220_),
    .B1(_03145_),
    .B2(_03147_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00125_));
 sky130_fd_sc_hd__a21oi_1 _08549_ (.A1(\sha256cu.K[30] ),
    .A2(_03139_),
    .B1(_03138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03148_));
 sky130_fd_sc_hd__a21oi_1 _08550_ (.A1(_03120_),
    .A2(_03122_),
    .B1(_03129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03149_));
 sky130_fd_sc_hd__o21a_1 _08551_ (.A1(_03134_),
    .A2(_03136_),
    .B1(_03132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03150_));
 sky130_fd_sc_hd__xnor2_1 _08552_ (.A(_03149_),
    .B(_03150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03151_));
 sky130_fd_sc_hd__and2b_1 _08553_ (.A_N(_03117_),
    .B(_03119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03152_));
 sky130_fd_sc_hd__a21oi_1 _08554_ (.A1(\sha256cu.m_out_digest.h_in[30] ),
    .A2(_03116_),
    .B1(_03152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03153_));
 sky130_fd_sc_hd__and2b_1 _08555_ (.A_N(_03125_),
    .B(_03126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03154_));
 sky130_fd_sc_hd__a21oi_1 _08556_ (.A1(\sha256cu.iter_processing.w[30] ),
    .A2(_03127_),
    .B1(_03154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03155_));
 sky130_fd_sc_hd__xnor2_4 _08557_ (.A(\sha256cu.m_out_digest.e_in[10] ),
    .B(\sha256cu.m_out_digest.e_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03156_));
 sky130_fd_sc_hd__xnor2_2 _08558_ (.A(\sha256cu.m_out_digest.e_in[24] ),
    .B(_03156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03157_));
 sky130_fd_sc_hd__mux2_1 _08559_ (.A0(\sha256cu.m_out_digest.g_in[31] ),
    .A1(\sha256cu.m_out_digest.f_in[31] ),
    .S(\sha256cu.m_out_digest.e_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03158_));
 sky130_fd_sc_hd__xnor2_1 _08560_ (.A(\sha256cu.iter_processing.w[31] ),
    .B(_03158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03159_));
 sky130_fd_sc_hd__xnor2_1 _08561_ (.A(_03157_),
    .B(_03159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03160_));
 sky130_fd_sc_hd__xnor2_1 _08562_ (.A(_03155_),
    .B(_03160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03161_));
 sky130_fd_sc_hd__xnor2_1 _08563_ (.A(_03153_),
    .B(_03161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03162_));
 sky130_fd_sc_hd__xor2_1 _08564_ (.A(_02382_),
    .B(\sha256cu.m_out_digest.a_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03163_));
 sky130_fd_sc_hd__a21o_1 _08565_ (.A1(\sha256cu.m_out_digest.b_in[31] ),
    .A2(\sha256cu.m_out_digest.a_in[31] ),
    .B1(\sha256cu.m_out_digest.c_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03164_));
 sky130_fd_sc_hd__o21a_1 _08566_ (.A1(\sha256cu.m_out_digest.b_in[31] ),
    .A2(\sha256cu.m_out_digest.a_in[31] ),
    .B1(_03164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03165_));
 sky130_fd_sc_hd__xor2_1 _08567_ (.A(\sha256cu.K[31] ),
    .B(\sha256cu.m_out_digest.h_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03166_));
 sky130_fd_sc_hd__xnor2_1 _08568_ (.A(\sha256cu.m_out_digest.a_in[21] ),
    .B(_03166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03167_));
 sky130_fd_sc_hd__xnor2_1 _08569_ (.A(_03165_),
    .B(_03167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03168_));
 sky130_fd_sc_hd__xnor2_1 _08570_ (.A(_03163_),
    .B(_03168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03169_));
 sky130_fd_sc_hd__xnor2_1 _08571_ (.A(_03162_),
    .B(_03169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03170_));
 sky130_fd_sc_hd__xnor2_1 _08572_ (.A(_03151_),
    .B(_03170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03171_));
 sky130_fd_sc_hd__xnor2_1 _08573_ (.A(_03148_),
    .B(_03171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03172_));
 sky130_fd_sc_hd__a21oi_1 _08574_ (.A1(_03142_),
    .A2(_03145_),
    .B1(_03172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03173_));
 sky130_fd_sc_hd__and3_1 _08575_ (.A(_03142_),
    .B(_03145_),
    .C(_03172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03174_));
 sky130_fd_sc_hd__or2_1 _08576_ (.A(\sha256cu.m_out_digest.a_in[31] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03175_));
 sky130_fd_sc_hd__o311a_1 _08577_ (.A1(_02040_),
    .A2(_03173_),
    .A3(_03174_),
    .B1(_03175_),
    .C1(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00126_));
 sky130_fd_sc_hd__o22a_1 _08578_ (.A1(\sha256cu.m_out_digest.b_in[0] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(\sha256cu.m_out_digest.a_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00127_));
 sky130_fd_sc_hd__a22o_1 _08579_ (.A1(\sha256cu.m_out_digest.b_in[1] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(\sha256cu.m_out_digest.a_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00128_));
 sky130_fd_sc_hd__o22a_1 _08580_ (.A1(\sha256cu.m_out_digest.b_in[2] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(\sha256cu.m_out_digest.a_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00129_));
 sky130_fd_sc_hd__a22o_1 _08581_ (.A1(\sha256cu.m_out_digest.b_in[3] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(\sha256cu.m_out_digest.a_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _08582_ (.A1(\sha256cu.m_out_digest.b_in[4] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(\sha256cu.m_out_digest.a_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _08583_ (.A1(\sha256cu.m_out_digest.b_in[5] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(\sha256cu.m_out_digest.a_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _08584_ (.A1(\sha256cu.m_out_digest.b_in[6] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(\sha256cu.m_out_digest.a_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00133_));
 sky130_fd_sc_hd__o22a_1 _08585_ (.A1(\sha256cu.m_out_digest.b_in[7] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(\sha256cu.m_out_digest.a_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00134_));
 sky130_fd_sc_hd__a22o_1 _08586_ (.A1(\sha256cu.m_out_digest.b_in[8] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(\sha256cu.m_out_digest.a_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00135_));
 sky130_fd_sc_hd__o22a_1 _08587_ (.A1(\sha256cu.m_out_digest.b_in[9] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(\sha256cu.m_out_digest.a_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00136_));
 sky130_fd_sc_hd__o22a_1 _08588_ (.A1(\sha256cu.m_out_digest.b_in[10] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(\sha256cu.m_out_digest.a_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00137_));
 sky130_fd_sc_hd__o22a_1 _08589_ (.A1(\sha256cu.m_out_digest.b_in[11] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(\sha256cu.m_out_digest.a_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00138_));
 sky130_fd_sc_hd__a22o_1 _08590_ (.A1(\sha256cu.m_out_digest.b_in[12] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(_02382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00139_));
 sky130_fd_sc_hd__o22a_1 _08591_ (.A1(\sha256cu.m_out_digest.b_in[13] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(_02027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00140_));
 sky130_fd_sc_hd__a22o_1 _08592_ (.A1(\sha256cu.m_out_digest.b_in[14] ),
    .A2(_03031_),
    .B1(_02114_),
    .B2(\sha256cu.m_out_digest.a_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00141_));
 sky130_fd_sc_hd__o22a_1 _08593_ (.A1(\sha256cu.m_out_digest.b_in[15] ),
    .A2(_02370_),
    .B1(_02110_),
    .B2(_02084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00142_));
 sky130_fd_sc_hd__buf_4 _08594_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03176_));
 sky130_fd_sc_hd__o22a_1 _08595_ (.A1(\sha256cu.m_out_digest.b_in[16] ),
    .A2(_02370_),
    .B1(_03176_),
    .B2(_02128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00143_));
 sky130_fd_sc_hd__buf_4 _08596_ (.A(_02369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03177_));
 sky130_fd_sc_hd__o22a_1 _08597_ (.A1(\sha256cu.m_out_digest.b_in[17] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(_02162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00144_));
 sky130_fd_sc_hd__o22a_1 _08598_ (.A1(\sha256cu.m_out_digest.b_in[18] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(_02198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00145_));
 sky130_fd_sc_hd__buf_6 _08599_ (.A(_02113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03178_));
 sky130_fd_sc_hd__a22o_1 _08600_ (.A1(\sha256cu.m_out_digest.b_in[19] ),
    .A2(_03031_),
    .B1(_03178_),
    .B2(_02233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00146_));
 sky130_fd_sc_hd__buf_6 _08601_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03179_));
 sky130_fd_sc_hd__a22o_1 _08602_ (.A1(\sha256cu.m_out_digest.b_in[20] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(_02273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00147_));
 sky130_fd_sc_hd__o22a_1 _08603_ (.A1(\sha256cu.m_out_digest.b_in[21] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(\sha256cu.m_out_digest.a_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00148_));
 sky130_fd_sc_hd__o22a_1 _08604_ (.A1(\sha256cu.m_out_digest.b_in[22] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(_02026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00149_));
 sky130_fd_sc_hd__a22o_1 _08605_ (.A1(\sha256cu.m_out_digest.b_in[23] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(\sha256cu.m_out_digest.a_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00150_));
 sky130_fd_sc_hd__o22a_1 _08606_ (.A1(\sha256cu.m_out_digest.b_in[24] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(_02083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00151_));
 sky130_fd_sc_hd__o22a_1 _08607_ (.A1(\sha256cu.m_out_digest.b_in[25] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(\sha256cu.m_out_digest.a_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00152_));
 sky130_fd_sc_hd__a22o_1 _08608_ (.A1(\sha256cu.m_out_digest.b_in[26] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(_02161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00153_));
 sky130_fd_sc_hd__o22a_1 _08609_ (.A1(\sha256cu.m_out_digest.b_in[27] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(\sha256cu.m_out_digest.a_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00154_));
 sky130_fd_sc_hd__o22a_1 _08610_ (.A1(\sha256cu.m_out_digest.b_in[28] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(_02232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00155_));
 sky130_fd_sc_hd__o22a_1 _08611_ (.A1(\sha256cu.m_out_digest.b_in[29] ),
    .A2(_03177_),
    .B1(_03176_),
    .B2(_02272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00156_));
 sky130_fd_sc_hd__a22o_1 _08612_ (.A1(\sha256cu.m_out_digest.b_in[30] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(_02304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00157_));
 sky130_fd_sc_hd__buf_4 _08613_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03180_));
 sky130_fd_sc_hd__o22a_1 _08614_ (.A1(\sha256cu.m_out_digest.b_in[31] ),
    .A2(_03177_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.a_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00158_));
 sky130_fd_sc_hd__a22o_1 _08615_ (.A1(\sha256cu.m_out_digest.c_in[0] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(\sha256cu.m_out_digest.b_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00159_));
 sky130_fd_sc_hd__buf_4 _08616_ (.A(_02369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03181_));
 sky130_fd_sc_hd__o22a_1 _08617_ (.A1(\sha256cu.m_out_digest.c_in[1] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00160_));
 sky130_fd_sc_hd__a22o_1 _08618_ (.A1(\sha256cu.m_out_digest.c_in[2] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(\sha256cu.m_out_digest.b_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00161_));
 sky130_fd_sc_hd__a22o_1 _08619_ (.A1(\sha256cu.m_out_digest.c_in[3] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(\sha256cu.m_out_digest.b_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00162_));
 sky130_fd_sc_hd__o22a_1 _08620_ (.A1(\sha256cu.m_out_digest.c_in[4] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00163_));
 sky130_fd_sc_hd__o22a_1 _08621_ (.A1(\sha256cu.m_out_digest.c_in[5] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00164_));
 sky130_fd_sc_hd__o22a_1 _08622_ (.A1(\sha256cu.m_out_digest.c_in[6] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00165_));
 sky130_fd_sc_hd__a22o_1 _08623_ (.A1(\sha256cu.m_out_digest.c_in[7] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(\sha256cu.m_out_digest.b_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00166_));
 sky130_fd_sc_hd__o22a_1 _08624_ (.A1(\sha256cu.m_out_digest.c_in[8] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00167_));
 sky130_fd_sc_hd__o22a_1 _08625_ (.A1(\sha256cu.m_out_digest.c_in[9] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00168_));
 sky130_fd_sc_hd__a22o_1 _08626_ (.A1(\sha256cu.m_out_digest.c_in[10] ),
    .A2(_03179_),
    .B1(_03178_),
    .B2(\sha256cu.m_out_digest.b_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00169_));
 sky130_fd_sc_hd__buf_4 _08627_ (.A(_02113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03182_));
 sky130_fd_sc_hd__a22o_1 _08628_ (.A1(\sha256cu.m_out_digest.c_in[11] ),
    .A2(_03179_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00170_));
 sky130_fd_sc_hd__o22a_1 _08629_ (.A1(\sha256cu.m_out_digest.c_in[12] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00171_));
 sky130_fd_sc_hd__o22a_1 _08630_ (.A1(\sha256cu.m_out_digest.c_in[13] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00172_));
 sky130_fd_sc_hd__o22a_1 _08631_ (.A1(\sha256cu.m_out_digest.c_in[14] ),
    .A2(_03181_),
    .B1(_03180_),
    .B2(\sha256cu.m_out_digest.b_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00173_));
 sky130_fd_sc_hd__buf_4 _08632_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03183_));
 sky130_fd_sc_hd__o22a_1 _08633_ (.A1(\sha256cu.m_out_digest.c_in[15] ),
    .A2(_03181_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00174_));
 sky130_fd_sc_hd__clkbuf_8 _08634_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03184_));
 sky130_fd_sc_hd__a22o_1 _08635_ (.A1(\sha256cu.m_out_digest.c_in[16] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00175_));
 sky130_fd_sc_hd__buf_4 _08636_ (.A(_02369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03185_));
 sky130_fd_sc_hd__o22a_1 _08637_ (.A1(\sha256cu.m_out_digest.c_in[17] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00176_));
 sky130_fd_sc_hd__o22a_1 _08638_ (.A1(\sha256cu.m_out_digest.c_in[18] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00177_));
 sky130_fd_sc_hd__o22a_1 _08639_ (.A1(\sha256cu.m_out_digest.c_in[19] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00178_));
 sky130_fd_sc_hd__a22o_1 _08640_ (.A1(\sha256cu.m_out_digest.c_in[20] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00179_));
 sky130_fd_sc_hd__o22a_1 _08641_ (.A1(\sha256cu.m_out_digest.c_in[21] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00180_));
 sky130_fd_sc_hd__o22a_1 _08642_ (.A1(\sha256cu.m_out_digest.c_in[22] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00181_));
 sky130_fd_sc_hd__a22o_1 _08643_ (.A1(\sha256cu.m_out_digest.c_in[23] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00182_));
 sky130_fd_sc_hd__a22o_1 _08644_ (.A1(\sha256cu.m_out_digest.c_in[24] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00183_));
 sky130_fd_sc_hd__a22o_1 _08645_ (.A1(\sha256cu.m_out_digest.c_in[25] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00184_));
 sky130_fd_sc_hd__o22a_1 _08646_ (.A1(\sha256cu.m_out_digest.c_in[26] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00185_));
 sky130_fd_sc_hd__o22a_1 _08647_ (.A1(\sha256cu.m_out_digest.c_in[27] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00186_));
 sky130_fd_sc_hd__o22a_1 _08648_ (.A1(\sha256cu.m_out_digest.c_in[28] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00187_));
 sky130_fd_sc_hd__o22a_1 _08649_ (.A1(\sha256cu.m_out_digest.c_in[29] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\sha256cu.m_out_digest.b_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00188_));
 sky130_fd_sc_hd__a22o_1 _08650_ (.A1(\sha256cu.m_out_digest.c_in[30] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00189_));
 sky130_fd_sc_hd__a22o_1 _08651_ (.A1(\sha256cu.m_out_digest.c_in[31] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.b_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00190_));
 sky130_fd_sc_hd__a22o_1 _08652_ (.A1(\sha256cu.m_out_digest.d_in[0] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.c_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00191_));
 sky130_fd_sc_hd__buf_4 _08653_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03186_));
 sky130_fd_sc_hd__o22a_1 _08654_ (.A1(\sha256cu.m_out_digest.d_in[1] ),
    .A2(_03185_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00192_));
 sky130_fd_sc_hd__a22o_1 _08655_ (.A1(\sha256cu.m_out_digest.d_in[2] ),
    .A2(_03184_),
    .B1(_03182_),
    .B2(\sha256cu.m_out_digest.c_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00193_));
 sky130_fd_sc_hd__buf_4 _08656_ (.A(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03187_));
 sky130_fd_sc_hd__o22a_1 _08657_ (.A1(\sha256cu.m_out_digest.d_in[3] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00194_));
 sky130_fd_sc_hd__o22a_1 _08658_ (.A1(\sha256cu.m_out_digest.d_in[4] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00195_));
 sky130_fd_sc_hd__o22a_1 _08659_ (.A1(\sha256cu.m_out_digest.d_in[5] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00196_));
 sky130_fd_sc_hd__buf_6 _08660_ (.A(_02113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03188_));
 sky130_fd_sc_hd__a22o_1 _08661_ (.A1(\sha256cu.m_out_digest.d_in[6] ),
    .A2(_03184_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00197_));
 sky130_fd_sc_hd__buf_6 _08662_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03189_));
 sky130_fd_sc_hd__a22o_1 _08663_ (.A1(\sha256cu.m_out_digest.d_in[7] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00198_));
 sky130_fd_sc_hd__o22a_1 _08664_ (.A1(\sha256cu.m_out_digest.d_in[8] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00199_));
 sky130_fd_sc_hd__a22o_1 _08665_ (.A1(\sha256cu.m_out_digest.d_in[9] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00200_));
 sky130_fd_sc_hd__o22a_1 _08666_ (.A1(\sha256cu.m_out_digest.d_in[10] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00201_));
 sky130_fd_sc_hd__a22o_1 _08667_ (.A1(\sha256cu.m_out_digest.d_in[11] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00202_));
 sky130_fd_sc_hd__o22a_1 _08668_ (.A1(\sha256cu.m_out_digest.d_in[12] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00203_));
 sky130_fd_sc_hd__o22a_1 _08669_ (.A1(\sha256cu.m_out_digest.d_in[13] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00204_));
 sky130_fd_sc_hd__o22a_1 _08670_ (.A1(\sha256cu.m_out_digest.d_in[14] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00205_));
 sky130_fd_sc_hd__o22a_1 _08671_ (.A1(\sha256cu.m_out_digest.d_in[15] ),
    .A2(_03187_),
    .B1(_03186_),
    .B2(\sha256cu.m_out_digest.c_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00206_));
 sky130_fd_sc_hd__buf_4 _08672_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03190_));
 sky130_fd_sc_hd__o22a_1 _08673_ (.A1(\sha256cu.m_out_digest.d_in[16] ),
    .A2(_03187_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00207_));
 sky130_fd_sc_hd__clkbuf_8 _08674_ (.A(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03191_));
 sky130_fd_sc_hd__o22a_1 _08675_ (.A1(\sha256cu.m_out_digest.d_in[17] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00208_));
 sky130_fd_sc_hd__o22a_1 _08676_ (.A1(\sha256cu.m_out_digest.d_in[18] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00209_));
 sky130_fd_sc_hd__o22a_1 _08677_ (.A1(\sha256cu.m_out_digest.d_in[19] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00210_));
 sky130_fd_sc_hd__a22o_1 _08678_ (.A1(\sha256cu.m_out_digest.d_in[20] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00211_));
 sky130_fd_sc_hd__a22o_1 _08679_ (.A1(\sha256cu.m_out_digest.d_in[21] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00212_));
 sky130_fd_sc_hd__o22a_1 _08680_ (.A1(\sha256cu.m_out_digest.d_in[22] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00213_));
 sky130_fd_sc_hd__a22o_1 _08681_ (.A1(\sha256cu.m_out_digest.d_in[23] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00214_));
 sky130_fd_sc_hd__o22a_1 _08682_ (.A1(\sha256cu.m_out_digest.d_in[24] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00215_));
 sky130_fd_sc_hd__a22o_1 _08683_ (.A1(\sha256cu.m_out_digest.d_in[25] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00216_));
 sky130_fd_sc_hd__o22a_1 _08684_ (.A1(\sha256cu.m_out_digest.d_in[26] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00217_));
 sky130_fd_sc_hd__a22o_1 _08685_ (.A1(\sha256cu.m_out_digest.d_in[27] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00218_));
 sky130_fd_sc_hd__a22o_1 _08686_ (.A1(\sha256cu.m_out_digest.d_in[28] ),
    .A2(_03189_),
    .B1(_03188_),
    .B2(\sha256cu.m_out_digest.c_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00219_));
 sky130_fd_sc_hd__o22a_1 _08687_ (.A1(\sha256cu.m_out_digest.d_in[29] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00220_));
 sky130_fd_sc_hd__buf_4 _08688_ (.A(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03192_));
 sky130_fd_sc_hd__a22o_1 _08689_ (.A1(\sha256cu.m_out_digest.d_in[30] ),
    .A2(_03189_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.c_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00221_));
 sky130_fd_sc_hd__o22a_1 _08690_ (.A1(\sha256cu.m_out_digest.d_in[31] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.c_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00222_));
 sky130_fd_sc_hd__nand2_1 _08691_ (.A(\sha256cu.iter_processing.w[0] ),
    .B(_02020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03193_));
 sky130_fd_sc_hd__or2_1 _08692_ (.A(\sha256cu.iter_processing.w[0] ),
    .B(_02020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03194_));
 sky130_fd_sc_hd__a21o_1 _08693_ (.A1(_03193_),
    .A2(_03194_),
    .B1(\sha256cu.K[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03195_));
 sky130_fd_sc_hd__nand3_1 _08694_ (.A(\sha256cu.K[0] ),
    .B(_03193_),
    .C(_03194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03196_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(_03195_),
    .B(_03196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03197_));
 sky130_fd_sc_hd__nand2_1 _08696_ (.A(\sha256cu.m_out_digest.h_in[0] ),
    .B(\sha256cu.m_out_digest.d_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03198_));
 sky130_fd_sc_hd__or2_1 _08697_ (.A(\sha256cu.m_out_digest.h_in[0] ),
    .B(\sha256cu.m_out_digest.d_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03199_));
 sky130_fd_sc_hd__nand2_1 _08698_ (.A(_03198_),
    .B(_03199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03200_));
 sky130_fd_sc_hd__xor2_1 _08699_ (.A(_02024_),
    .B(_03200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03201_));
 sky130_fd_sc_hd__nor2_1 _08700_ (.A(_03197_),
    .B(_03201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03202_));
 sky130_fd_sc_hd__a21o_1 _08701_ (.A1(_03197_),
    .A2(_03201_),
    .B1(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03203_));
 sky130_fd_sc_hd__a21oi_1 _08702_ (.A1(\sha256cu.m_out_digest.e_in[0] ),
    .A2(_02732_),
    .B1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03204_));
 sky130_fd_sc_hd__o21ai_1 _08703_ (.A1(_03202_),
    .A2(_03203_),
    .B1(_03204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00223_));
 sky130_fd_sc_hd__nand2_1 _08704_ (.A(\sha256cu.m_out_digest.h_in[1] ),
    .B(\sha256cu.m_out_digest.d_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03205_));
 sky130_fd_sc_hd__or2_1 _08705_ (.A(\sha256cu.m_out_digest.h_in[1] ),
    .B(\sha256cu.m_out_digest.d_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03206_));
 sky130_fd_sc_hd__nand2_1 _08706_ (.A(_03205_),
    .B(_03206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03207_));
 sky130_fd_sc_hd__xor2_1 _08707_ (.A(_02051_),
    .B(_03207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03208_));
 sky130_fd_sc_hd__a21boi_1 _08708_ (.A1(_02024_),
    .A2(_03199_),
    .B1_N(_03198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03209_));
 sky130_fd_sc_hd__xnor2_1 _08709_ (.A(_03208_),
    .B(_03209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03210_));
 sky130_fd_sc_hd__inv_2 _08710_ (.A(\sha256cu.K[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03211_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(\sha256cu.iter_processing.w[1] ),
    .B(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03212_));
 sky130_fd_sc_hd__or2_1 _08712_ (.A(\sha256cu.iter_processing.w[1] ),
    .B(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03213_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(_03212_),
    .B(_03213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03214_));
 sky130_fd_sc_hd__xnor2_1 _08714_ (.A(_03211_),
    .B(_03214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03215_));
 sky130_fd_sc_hd__xor2_1 _08715_ (.A(_03210_),
    .B(_03215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03216_));
 sky130_fd_sc_hd__xnor2_1 _08716_ (.A(_03202_),
    .B(_03216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03217_));
 sky130_fd_sc_hd__a21o_1 _08717_ (.A1(_03193_),
    .A2(_03196_),
    .B1(_03217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03218_));
 sky130_fd_sc_hd__a31oi_1 _08718_ (.A1(_03193_),
    .A2(_03196_),
    .A3(_03217_),
    .B1(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03219_));
 sky130_fd_sc_hd__a221o_1 _08719_ (.A1(\sha256cu.m_out_digest.e_in[1] ),
    .A2(_02220_),
    .B1(_03218_),
    .B2(_03219_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00224_));
 sky130_fd_sc_hd__nand2_1 _08720_ (.A(_03202_),
    .B(_03216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03220_));
 sky130_fd_sc_hd__o21ai_1 _08721_ (.A1(_03211_),
    .A2(_03214_),
    .B1(_03212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03221_));
 sky130_fd_sc_hd__nand2_1 _08722_ (.A(\sha256cu.iter_processing.w[2] ),
    .B(_02075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03222_));
 sky130_fd_sc_hd__or2_1 _08723_ (.A(\sha256cu.iter_processing.w[2] ),
    .B(_02075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03223_));
 sky130_fd_sc_hd__nand2_1 _08724_ (.A(_03222_),
    .B(_03223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03224_));
 sky130_fd_sc_hd__xnor2_1 _08725_ (.A(_02071_),
    .B(_03224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03225_));
 sky130_fd_sc_hd__nand2_1 _08726_ (.A(\sha256cu.m_out_digest.h_in[2] ),
    .B(\sha256cu.m_out_digest.d_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03226_));
 sky130_fd_sc_hd__or2_1 _08727_ (.A(\sha256cu.m_out_digest.h_in[2] ),
    .B(\sha256cu.m_out_digest.d_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03227_));
 sky130_fd_sc_hd__nand2_1 _08728_ (.A(_03226_),
    .B(_03227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03228_));
 sky130_fd_sc_hd__xor2_1 _08729_ (.A(_02081_),
    .B(_03228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03229_));
 sky130_fd_sc_hd__a21boi_1 _08730_ (.A1(_02051_),
    .A2(_03206_),
    .B1_N(_03205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03230_));
 sky130_fd_sc_hd__xnor2_1 _08731_ (.A(_03229_),
    .B(_03230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03231_));
 sky130_fd_sc_hd__xor2_1 _08732_ (.A(_03225_),
    .B(_03231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03232_));
 sky130_fd_sc_hd__or2_1 _08733_ (.A(_03208_),
    .B(_03209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03233_));
 sky130_fd_sc_hd__o21ai_1 _08734_ (.A1(_03210_),
    .A2(_03215_),
    .B1(_03233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03234_));
 sky130_fd_sc_hd__xor2_1 _08735_ (.A(_03232_),
    .B(_03234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03235_));
 sky130_fd_sc_hd__xnor2_1 _08736_ (.A(_03221_),
    .B(_03235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03236_));
 sky130_fd_sc_hd__a21oi_2 _08737_ (.A1(_03220_),
    .A2(_03218_),
    .B1(_03236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03237_));
 sky130_fd_sc_hd__a31o_1 _08738_ (.A1(_03220_),
    .A2(_03218_),
    .A3(_03236_),
    .B1(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03238_));
 sky130_fd_sc_hd__nor2_1 _08739_ (.A(_03237_),
    .B(_03238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03239_));
 sky130_fd_sc_hd__a211o_1 _08740_ (.A1(\sha256cu.m_out_digest.e_in[2] ),
    .A2(_02040_),
    .B1(_03239_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00225_));
 sky130_fd_sc_hd__o21ai_2 _08741_ (.A1(_02071_),
    .A2(_03224_),
    .B1(_03222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03240_));
 sky130_fd_sc_hd__nand2_1 _08742_ (.A(\sha256cu.iter_processing.w[3] ),
    .B(_02120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03241_));
 sky130_fd_sc_hd__or2_1 _08743_ (.A(\sha256cu.iter_processing.w[3] ),
    .B(_02120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03242_));
 sky130_fd_sc_hd__nand2_1 _08744_ (.A(_03241_),
    .B(_03242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03243_));
 sky130_fd_sc_hd__xor2_1 _08745_ (.A(\sha256cu.K[3] ),
    .B(_03243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03244_));
 sky130_fd_sc_hd__or2_1 _08746_ (.A(\sha256cu.m_out_digest.h_in[3] ),
    .B(\sha256cu.m_out_digest.d_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03245_));
 sky130_fd_sc_hd__nand2_1 _08747_ (.A(\sha256cu.m_out_digest.h_in[3] ),
    .B(\sha256cu.m_out_digest.d_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03246_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(_03245_),
    .B(_03246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03247_));
 sky130_fd_sc_hd__xor2_1 _08749_ (.A(_02126_),
    .B(_03247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03248_));
 sky130_fd_sc_hd__a21boi_1 _08750_ (.A1(_02081_),
    .A2(_03227_),
    .B1_N(_03226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03249_));
 sky130_fd_sc_hd__xnor2_1 _08751_ (.A(_03248_),
    .B(_03249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03250_));
 sky130_fd_sc_hd__xor2_1 _08752_ (.A(_03244_),
    .B(_03250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03251_));
 sky130_fd_sc_hd__or2_1 _08753_ (.A(_03229_),
    .B(_03230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03252_));
 sky130_fd_sc_hd__o21a_1 _08754_ (.A1(_03225_),
    .A2(_03231_),
    .B1(_03252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03253_));
 sky130_fd_sc_hd__xnor2_1 _08755_ (.A(_03251_),
    .B(_03253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03254_));
 sky130_fd_sc_hd__xnor2_1 _08756_ (.A(_03240_),
    .B(_03254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03255_));
 sky130_fd_sc_hd__nand2_1 _08757_ (.A(_03232_),
    .B(_03234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03256_));
 sky130_fd_sc_hd__a21boi_1 _08758_ (.A1(_03221_),
    .A2(_03235_),
    .B1_N(_03256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03257_));
 sky130_fd_sc_hd__xor2_1 _08759_ (.A(_03255_),
    .B(_03257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03258_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_03237_),
    .B(_03258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03259_));
 sky130_fd_sc_hd__o21a_1 _08761_ (.A1(_03237_),
    .A2(_03258_),
    .B1(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03260_));
 sky130_fd_sc_hd__a221o_1 _08762_ (.A1(\sha256cu.m_out_digest.e_in[3] ),
    .A2(_02732_),
    .B1(_03259_),
    .B2(_03260_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00226_));
 sky130_fd_sc_hd__inv_2 _08763_ (.A(\sha256cu.m_out_digest.e_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03261_));
 sky130_fd_sc_hd__nor2_1 _08764_ (.A(_03255_),
    .B(_03257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03262_));
 sky130_fd_sc_hd__a21o_1 _08765_ (.A1(_03237_),
    .A2(_03258_),
    .B1(_03262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03263_));
 sky130_fd_sc_hd__a21bo_1 _08766_ (.A1(\sha256cu.K[3] ),
    .A2(_03242_),
    .B1_N(_03241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03264_));
 sky130_fd_sc_hd__or2_1 _08767_ (.A(\sha256cu.m_out_digest.h_in[4] ),
    .B(\sha256cu.m_out_digest.d_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03265_));
 sky130_fd_sc_hd__nand2_1 _08768_ (.A(\sha256cu.m_out_digest.h_in[4] ),
    .B(\sha256cu.m_out_digest.d_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _08769_ (.A(_03265_),
    .B(_03266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03267_));
 sky130_fd_sc_hd__xor2_1 _08770_ (.A(_02159_),
    .B(_03267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03268_));
 sky130_fd_sc_hd__a21boi_1 _08771_ (.A1(_02126_),
    .A2(_03245_),
    .B1_N(_03246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03269_));
 sky130_fd_sc_hd__xnor2_1 _08772_ (.A(_03268_),
    .B(_03269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03270_));
 sky130_fd_sc_hd__inv_2 _08773_ (.A(\sha256cu.K[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03271_));
 sky130_fd_sc_hd__or2_1 _08774_ (.A(\sha256cu.iter_processing.w[4] ),
    .B(_02153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03272_));
 sky130_fd_sc_hd__nand2_1 _08775_ (.A(\sha256cu.iter_processing.w[4] ),
    .B(_02153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03273_));
 sky130_fd_sc_hd__nand2_1 _08776_ (.A(_03272_),
    .B(_03273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03274_));
 sky130_fd_sc_hd__xnor2_1 _08777_ (.A(_03271_),
    .B(_03274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03275_));
 sky130_fd_sc_hd__xor2_1 _08778_ (.A(_03270_),
    .B(_03275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03276_));
 sky130_fd_sc_hd__or2_1 _08779_ (.A(_03248_),
    .B(_03249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03277_));
 sky130_fd_sc_hd__o21a_1 _08780_ (.A1(_03244_),
    .A2(_03250_),
    .B1(_03277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03278_));
 sky130_fd_sc_hd__xnor2_1 _08781_ (.A(_03276_),
    .B(_03278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03279_));
 sky130_fd_sc_hd__nand2_1 _08782_ (.A(_03264_),
    .B(_03279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03280_));
 sky130_fd_sc_hd__or2_1 _08783_ (.A(_03264_),
    .B(_03279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03281_));
 sky130_fd_sc_hd__nand2_1 _08784_ (.A(_03280_),
    .B(_03281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03282_));
 sky130_fd_sc_hd__or2b_1 _08785_ (.A(_03253_),
    .B_N(_03251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03283_));
 sky130_fd_sc_hd__a21boi_2 _08786_ (.A1(_03240_),
    .A2(_03254_),
    .B1_N(_03283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03284_));
 sky130_fd_sc_hd__xor2_2 _08787_ (.A(_03282_),
    .B(_03284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03285_));
 sky130_fd_sc_hd__and2_1 _08788_ (.A(_03263_),
    .B(_03285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03286_));
 sky130_fd_sc_hd__o21ai_1 _08789_ (.A1(_03263_),
    .A2(_03285_),
    .B1(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03287_));
 sky130_fd_sc_hd__buf_4 _08790_ (.A(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03288_));
 sky130_fd_sc_hd__o221a_1 _08791_ (.A1(_03261_),
    .A2(_02440_),
    .B1(_03286_),
    .B2(_03287_),
    .C1(_03288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03289_));
 sky130_fd_sc_hd__inv_1 _08792_ (.A(_03289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00227_));
 sky130_fd_sc_hd__or2b_1 _08793_ (.A(_03278_),
    .B_N(_03276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03290_));
 sky130_fd_sc_hd__nor2_1 _08794_ (.A(\sha256cu.m_out_digest.h_in[5] ),
    .B(\sha256cu.m_out_digest.d_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03291_));
 sky130_fd_sc_hd__and2_1 _08795_ (.A(\sha256cu.m_out_digest.h_in[5] ),
    .B(\sha256cu.m_out_digest.d_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03292_));
 sky130_fd_sc_hd__nor2_1 _08796_ (.A(_03291_),
    .B(_03292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03293_));
 sky130_fd_sc_hd__xnor2_1 _08797_ (.A(_02196_),
    .B(_03293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03294_));
 sky130_fd_sc_hd__a21boi_1 _08798_ (.A1(_02159_),
    .A2(_03265_),
    .B1_N(_03266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03295_));
 sky130_fd_sc_hd__xnor2_1 _08799_ (.A(_03294_),
    .B(_03295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03296_));
 sky130_fd_sc_hd__and2_1 _08800_ (.A(\sha256cu.iter_processing.w[5] ),
    .B(_02190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03297_));
 sky130_fd_sc_hd__or2_1 _08801_ (.A(\sha256cu.iter_processing.w[5] ),
    .B(_02190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03298_));
 sky130_fd_sc_hd__or2b_1 _08802_ (.A(_03297_),
    .B_N(_03298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03299_));
 sky130_fd_sc_hd__xor2_1 _08803_ (.A(\sha256cu.K[5] ),
    .B(_03299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03300_));
 sky130_fd_sc_hd__xor2_1 _08804_ (.A(_03296_),
    .B(_03300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03301_));
 sky130_fd_sc_hd__or2_1 _08805_ (.A(_03268_),
    .B(_03269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03302_));
 sky130_fd_sc_hd__o21a_1 _08806_ (.A1(_03270_),
    .A2(_03275_),
    .B1(_03302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03303_));
 sky130_fd_sc_hd__xnor2_1 _08807_ (.A(_03301_),
    .B(_03303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03304_));
 sky130_fd_sc_hd__o21ai_1 _08808_ (.A1(_03271_),
    .A2(_03274_),
    .B1(_03273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03305_));
 sky130_fd_sc_hd__xnor2_1 _08809_ (.A(_03304_),
    .B(_03305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03306_));
 sky130_fd_sc_hd__a21oi_2 _08810_ (.A1(_03290_),
    .A2(_03280_),
    .B1(_03306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03307_));
 sky130_fd_sc_hd__and3_1 _08811_ (.A(_03290_),
    .B(_03280_),
    .C(_03306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03308_));
 sky130_fd_sc_hd__nor2_1 _08812_ (.A(_03307_),
    .B(_03308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03309_));
 sky130_fd_sc_hd__o21ba_1 _08813_ (.A1(_03282_),
    .A2(_03284_),
    .B1_N(_03286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03310_));
 sky130_fd_sc_hd__xnor2_1 _08814_ (.A(_03309_),
    .B(_03310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03311_));
 sky130_fd_sc_hd__a22o_1 _08815_ (.A1(\sha256cu.m_out_digest.e_in[5] ),
    .A2(_02037_),
    .B1(_02017_),
    .B2(_03311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03312_));
 sky130_fd_sc_hd__or2_1 _08816_ (.A(_02002_),
    .B(_03312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_1 _08817_ (.A(_03313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00228_));
 sky130_fd_sc_hd__nor3_1 _08818_ (.A(_03282_),
    .B(_03284_),
    .C(_03308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03314_));
 sky130_fd_sc_hd__a311oi_4 _08819_ (.A1(_03263_),
    .A2(_03285_),
    .A3(_03309_),
    .B1(_03314_),
    .C1(_03307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03315_));
 sky130_fd_sc_hd__nor2_1 _08820_ (.A(_03294_),
    .B(_03295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03316_));
 sky130_fd_sc_hd__nor2_1 _08821_ (.A(_03296_),
    .B(_03300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03317_));
 sky130_fd_sc_hd__nor2_1 _08822_ (.A(\sha256cu.iter_processing.w[6] ),
    .B(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03318_));
 sky130_fd_sc_hd__and2_1 _08823_ (.A(\sha256cu.iter_processing.w[6] ),
    .B(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03319_));
 sky130_fd_sc_hd__nor2_1 _08824_ (.A(_03318_),
    .B(_03319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03320_));
 sky130_fd_sc_hd__xnor2_1 _08825_ (.A(\sha256cu.K[6] ),
    .B(_03320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03321_));
 sky130_fd_sc_hd__nor2_1 _08826_ (.A(\sha256cu.m_out_digest.h_in[6] ),
    .B(\sha256cu.m_out_digest.d_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03322_));
 sky130_fd_sc_hd__and2_1 _08827_ (.A(\sha256cu.m_out_digest.h_in[6] ),
    .B(\sha256cu.m_out_digest.d_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03323_));
 sky130_fd_sc_hd__nor2_1 _08828_ (.A(_03322_),
    .B(_03323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03324_));
 sky130_fd_sc_hd__xnor2_1 _08829_ (.A(_02230_),
    .B(_03324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03325_));
 sky130_fd_sc_hd__a21oi_1 _08830_ (.A1(_02196_),
    .A2(_03293_),
    .B1(_03292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03326_));
 sky130_fd_sc_hd__xnor2_1 _08831_ (.A(_03325_),
    .B(_03326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03327_));
 sky130_fd_sc_hd__xor2_1 _08832_ (.A(_03321_),
    .B(_03327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03328_));
 sky130_fd_sc_hd__o21ai_1 _08833_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03329_));
 sky130_fd_sc_hd__or3_1 _08834_ (.A(_03316_),
    .B(_03317_),
    .C(_03328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03330_));
 sky130_fd_sc_hd__and2_1 _08835_ (.A(_03329_),
    .B(_03330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03331_));
 sky130_fd_sc_hd__a21o_1 _08836_ (.A1(\sha256cu.K[5] ),
    .A2(_03298_),
    .B1(_03297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03332_));
 sky130_fd_sc_hd__xor2_1 _08837_ (.A(_03331_),
    .B(_03332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03333_));
 sky130_fd_sc_hd__or2b_1 _08838_ (.A(_03303_),
    .B_N(_03301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03334_));
 sky130_fd_sc_hd__a21bo_1 _08839_ (.A1(_03304_),
    .A2(_03305_),
    .B1_N(_03334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03335_));
 sky130_fd_sc_hd__nand2_1 _08840_ (.A(_03333_),
    .B(_03335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03336_));
 sky130_fd_sc_hd__or2_1 _08841_ (.A(_03333_),
    .B(_03335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03337_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(_03336_),
    .B(_03337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03338_));
 sky130_fd_sc_hd__or2_1 _08843_ (.A(_03315_),
    .B(_03338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03339_));
 sky130_fd_sc_hd__a21oi_1 _08844_ (.A1(_03315_),
    .A2(_03338_),
    .B1(_02732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03340_));
 sky130_fd_sc_hd__a221o_1 _08845_ (.A1(\sha256cu.m_out_digest.e_in[6] ),
    .A2(_02732_),
    .B1(_03339_),
    .B2(_03340_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00229_));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(_03331_),
    .B(_03332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03341_));
 sky130_fd_sc_hd__a21o_1 _08847_ (.A1(\sha256cu.K[6] ),
    .A2(_03320_),
    .B1(_03319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03342_));
 sky130_fd_sc_hd__nor2_1 _08848_ (.A(_03325_),
    .B(_03326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03343_));
 sky130_fd_sc_hd__nor2_1 _08849_ (.A(_03321_),
    .B(_03327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03344_));
 sky130_fd_sc_hd__nand2_1 _08850_ (.A(\sha256cu.iter_processing.w[7] ),
    .B(_02264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03345_));
 sky130_fd_sc_hd__or2_1 _08851_ (.A(\sha256cu.iter_processing.w[7] ),
    .B(_02264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03346_));
 sky130_fd_sc_hd__nand2_1 _08852_ (.A(_03345_),
    .B(_03346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03347_));
 sky130_fd_sc_hd__xor2_1 _08853_ (.A(\sha256cu.K[7] ),
    .B(_03347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03348_));
 sky130_fd_sc_hd__or2_1 _08854_ (.A(\sha256cu.m_out_digest.h_in[7] ),
    .B(\sha256cu.m_out_digest.d_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03349_));
 sky130_fd_sc_hd__nand2_1 _08855_ (.A(\sha256cu.m_out_digest.h_in[7] ),
    .B(\sha256cu.m_out_digest.d_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03350_));
 sky130_fd_sc_hd__nand2_1 _08856_ (.A(_03349_),
    .B(_03350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03351_));
 sky130_fd_sc_hd__xor2_1 _08857_ (.A(_02270_),
    .B(_03351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03352_));
 sky130_fd_sc_hd__a21oi_1 _08858_ (.A1(_02230_),
    .A2(_03324_),
    .B1(_03323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03353_));
 sky130_fd_sc_hd__xnor2_1 _08859_ (.A(_03352_),
    .B(_03353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03354_));
 sky130_fd_sc_hd__xor2_1 _08860_ (.A(_03348_),
    .B(_03354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03355_));
 sky130_fd_sc_hd__o21ai_1 _08861_ (.A1(_03343_),
    .A2(_03344_),
    .B1(_03355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03356_));
 sky130_fd_sc_hd__or3_1 _08862_ (.A(_03343_),
    .B(_03344_),
    .C(_03355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03357_));
 sky130_fd_sc_hd__and2_1 _08863_ (.A(_03356_),
    .B(_03357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03358_));
 sky130_fd_sc_hd__xnor2_1 _08864_ (.A(_03342_),
    .B(_03358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03359_));
 sky130_fd_sc_hd__and3_1 _08865_ (.A(_03329_),
    .B(_03341_),
    .C(_03359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03360_));
 sky130_fd_sc_hd__a21o_1 _08866_ (.A1(_03329_),
    .A2(_03341_),
    .B1(_03359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03361_));
 sky130_fd_sc_hd__or2b_1 _08867_ (.A(_03360_),
    .B_N(_03361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03362_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(_03336_),
    .B(_03339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03363_));
 sky130_fd_sc_hd__xnor2_1 _08869_ (.A(_03362_),
    .B(_03363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03364_));
 sky130_fd_sc_hd__or2_1 _08870_ (.A(\sha256cu.m_out_digest.e_in[7] ),
    .B(_02440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_8 _08871_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03366_));
 sky130_fd_sc_hd__o211a_1 _08872_ (.A1(_02332_),
    .A2(_03364_),
    .B1(_03365_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00230_));
 sky130_fd_sc_hd__nand2_1 _08873_ (.A(_03342_),
    .B(_03358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03367_));
 sky130_fd_sc_hd__a21bo_1 _08874_ (.A1(\sha256cu.K[7] ),
    .A2(_03346_),
    .B1_N(_03345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03368_));
 sky130_fd_sc_hd__or2_1 _08875_ (.A(\sha256cu.m_out_digest.h_in[8] ),
    .B(\sha256cu.m_out_digest.d_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03369_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(\sha256cu.m_out_digest.h_in[8] ),
    .B(\sha256cu.m_out_digest.d_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03370_));
 sky130_fd_sc_hd__nand2_1 _08877_ (.A(_03369_),
    .B(_03370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03371_));
 sky130_fd_sc_hd__xor2_1 _08878_ (.A(_02302_),
    .B(_03371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03372_));
 sky130_fd_sc_hd__a21bo_1 _08879_ (.A1(_02270_),
    .A2(_03349_),
    .B1_N(_03350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03373_));
 sky130_fd_sc_hd__and2b_1 _08880_ (.A_N(_03372_),
    .B(_03373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03374_));
 sky130_fd_sc_hd__and2b_1 _08881_ (.A_N(_03373_),
    .B(_03372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03375_));
 sky130_fd_sc_hd__or2_1 _08882_ (.A(_03374_),
    .B(_03375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03376_));
 sky130_fd_sc_hd__inv_2 _08883_ (.A(\sha256cu.K[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _08884_ (.A(\sha256cu.iter_processing.w[8] ),
    .B(_02296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03378_));
 sky130_fd_sc_hd__or2_1 _08885_ (.A(\sha256cu.iter_processing.w[8] ),
    .B(_02296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03379_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(_03378_),
    .B(_03379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03380_));
 sky130_fd_sc_hd__xnor2_1 _08887_ (.A(_03377_),
    .B(_03380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03381_));
 sky130_fd_sc_hd__xor2_1 _08888_ (.A(_03376_),
    .B(_03381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03382_));
 sky130_fd_sc_hd__or2_1 _08889_ (.A(_03352_),
    .B(_03353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03383_));
 sky130_fd_sc_hd__o21a_1 _08890_ (.A1(_03348_),
    .A2(_03354_),
    .B1(_03383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03384_));
 sky130_fd_sc_hd__xnor2_1 _08891_ (.A(_03382_),
    .B(_03384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03385_));
 sky130_fd_sc_hd__xnor2_1 _08892_ (.A(_03368_),
    .B(_03385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03386_));
 sky130_fd_sc_hd__a21oi_1 _08893_ (.A1(_03356_),
    .A2(_03367_),
    .B1(_03386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03387_));
 sky130_fd_sc_hd__and3_1 _08894_ (.A(_03356_),
    .B(_03367_),
    .C(_03386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03388_));
 sky130_fd_sc_hd__nor2_1 _08895_ (.A(_03387_),
    .B(_03388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03389_));
 sky130_fd_sc_hd__a21o_1 _08896_ (.A1(_03336_),
    .A2(_03361_),
    .B1(_03360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03390_));
 sky130_fd_sc_hd__o31a_2 _08897_ (.A1(_03315_),
    .A2(_03338_),
    .A3(_03362_),
    .B1(_03390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03391_));
 sky130_fd_sc_hd__xnor2_1 _08898_ (.A(_03389_),
    .B(_03391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03392_));
 sky130_fd_sc_hd__or2_1 _08899_ (.A(\sha256cu.m_out_digest.e_in[8] ),
    .B(_02440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03393_));
 sky130_fd_sc_hd__o211a_1 _08900_ (.A1(_02040_),
    .A2(_03392_),
    .B1(_03393_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00231_));
 sky130_fd_sc_hd__or2b_1 _08901_ (.A(_03384_),
    .B_N(_03382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03394_));
 sky130_fd_sc_hd__nand2_1 _08902_ (.A(_03368_),
    .B(_03385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03395_));
 sky130_fd_sc_hd__or2_1 _08903_ (.A(\sha256cu.m_out_digest.h_in[9] ),
    .B(\sha256cu.m_out_digest.d_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03396_));
 sky130_fd_sc_hd__nand2_1 _08904_ (.A(\sha256cu.m_out_digest.h_in[9] ),
    .B(\sha256cu.m_out_digest.d_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _08905_ (.A(_03396_),
    .B(_03397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03398_));
 sky130_fd_sc_hd__xor2_1 _08906_ (.A(_02344_),
    .B(_03398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03399_));
 sky130_fd_sc_hd__a21boi_1 _08907_ (.A1(_02302_),
    .A2(_03369_),
    .B1_N(_03370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03400_));
 sky130_fd_sc_hd__nor2_1 _08908_ (.A(_03399_),
    .B(_03400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03401_));
 sky130_fd_sc_hd__nand2_1 _08909_ (.A(_03399_),
    .B(_03400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03402_));
 sky130_fd_sc_hd__or2b_1 _08910_ (.A(_03401_),
    .B_N(_03402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03403_));
 sky130_fd_sc_hd__or2_1 _08911_ (.A(\sha256cu.iter_processing.w[9] ),
    .B(_02338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03404_));
 sky130_fd_sc_hd__nand2_1 _08912_ (.A(\sha256cu.iter_processing.w[9] ),
    .B(_02338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _08913_ (.A(_03404_),
    .B(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03406_));
 sky130_fd_sc_hd__xor2_1 _08914_ (.A(\sha256cu.K[9] ),
    .B(_03406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03407_));
 sky130_fd_sc_hd__xor2_1 _08915_ (.A(_03403_),
    .B(_03407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03408_));
 sky130_fd_sc_hd__o21ba_1 _08916_ (.A1(_03375_),
    .A2(_03381_),
    .B1_N(_03374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03409_));
 sky130_fd_sc_hd__xnor2_1 _08917_ (.A(_03408_),
    .B(_03409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03410_));
 sky130_fd_sc_hd__o21ai_1 _08918_ (.A1(_03377_),
    .A2(_03380_),
    .B1(_03378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03411_));
 sky130_fd_sc_hd__xnor2_1 _08919_ (.A(_03410_),
    .B(_03411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03412_));
 sky130_fd_sc_hd__a21oi_1 _08920_ (.A1(_03394_),
    .A2(_03395_),
    .B1(_03412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03413_));
 sky130_fd_sc_hd__and3_1 _08921_ (.A(_03394_),
    .B(_03395_),
    .C(_03412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03414_));
 sky130_fd_sc_hd__nor2_1 _08922_ (.A(_03413_),
    .B(_03414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03415_));
 sky130_fd_sc_hd__a21o_1 _08923_ (.A1(_03356_),
    .A2(_03367_),
    .B1(_03386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03416_));
 sky130_fd_sc_hd__o21a_1 _08924_ (.A1(_03388_),
    .A2(_03391_),
    .B1(_03416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03417_));
 sky130_fd_sc_hd__xnor2_1 _08925_ (.A(_03415_),
    .B(_03417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03418_));
 sky130_fd_sc_hd__a22o_1 _08926_ (.A1(\sha256cu.m_out_digest.e_in[9] ),
    .A2(_02037_),
    .B1(_02017_),
    .B2(_03418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03419_));
 sky130_fd_sc_hd__or2_1 _08927_ (.A(_02002_),
    .B(_03419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_1 _08928_ (.A(_03420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00232_));
 sky130_fd_sc_hd__or2b_1 _08929_ (.A(_03409_),
    .B_N(_03408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03421_));
 sky130_fd_sc_hd__nand2_1 _08930_ (.A(_03410_),
    .B(_03411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03422_));
 sky130_fd_sc_hd__or2_1 _08931_ (.A(\sha256cu.m_out_digest.h_in[10] ),
    .B(\sha256cu.m_out_digest.d_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03423_));
 sky130_fd_sc_hd__nand2_1 _08932_ (.A(\sha256cu.m_out_digest.h_in[10] ),
    .B(\sha256cu.m_out_digest.d_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03424_));
 sky130_fd_sc_hd__nand2_1 _08933_ (.A(_03423_),
    .B(_03424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03425_));
 sky130_fd_sc_hd__xor2_1 _08934_ (.A(_02380_),
    .B(_03425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03426_));
 sky130_fd_sc_hd__a21boi_1 _08935_ (.A1(_02344_),
    .A2(_03396_),
    .B1_N(_03397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03427_));
 sky130_fd_sc_hd__nor2_1 _08936_ (.A(_03426_),
    .B(_03427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03428_));
 sky130_fd_sc_hd__nand2_1 _08937_ (.A(_03426_),
    .B(_03427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03429_));
 sky130_fd_sc_hd__or2b_1 _08938_ (.A(_03428_),
    .B_N(_03429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03430_));
 sky130_fd_sc_hd__inv_2 _08939_ (.A(\sha256cu.K[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03431_));
 sky130_fd_sc_hd__or2_1 _08940_ (.A(\sha256cu.iter_processing.w[10] ),
    .B(_02374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03432_));
 sky130_fd_sc_hd__nand2_1 _08941_ (.A(\sha256cu.iter_processing.w[10] ),
    .B(_02374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_1 _08942_ (.A(_03432_),
    .B(_03433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03434_));
 sky130_fd_sc_hd__xnor2_2 _08943_ (.A(_03431_),
    .B(_03434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03435_));
 sky130_fd_sc_hd__xor2_2 _08944_ (.A(_03430_),
    .B(_03435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03436_));
 sky130_fd_sc_hd__o21ba_1 _08945_ (.A1(_03403_),
    .A2(_03407_),
    .B1_N(_03401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03437_));
 sky130_fd_sc_hd__xnor2_1 _08946_ (.A(_03436_),
    .B(_03437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03438_));
 sky130_fd_sc_hd__a21bo_1 _08947_ (.A1(\sha256cu.K[9] ),
    .A2(_03404_),
    .B1_N(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03439_));
 sky130_fd_sc_hd__xnor2_1 _08948_ (.A(_03438_),
    .B(_03439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03440_));
 sky130_fd_sc_hd__a21o_1 _08949_ (.A1(_03421_),
    .A2(_03422_),
    .B1(_03440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03441_));
 sky130_fd_sc_hd__nand3_1 _08950_ (.A(_03421_),
    .B(_03422_),
    .C(_03440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03442_));
 sky130_fd_sc_hd__and2_1 _08951_ (.A(_03441_),
    .B(_03442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03443_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(_03389_),
    .B(_03415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03444_));
 sky130_fd_sc_hd__nor2_1 _08953_ (.A(_03391_),
    .B(_03444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03445_));
 sky130_fd_sc_hd__a21o_1 _08954_ (.A1(_03394_),
    .A2(_03395_),
    .B1(_03412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03446_));
 sky130_fd_sc_hd__a21oi_2 _08955_ (.A1(_03416_),
    .A2(_03446_),
    .B1(_03414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03447_));
 sky130_fd_sc_hd__o21ai_1 _08956_ (.A1(_03445_),
    .A2(_03447_),
    .B1(_03443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03448_));
 sky130_fd_sc_hd__o311a_1 _08957_ (.A1(_03443_),
    .A2(_03445_),
    .A3(_03447_),
    .B1(_03448_),
    .C1(_02113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03449_));
 sky130_fd_sc_hd__a21o_1 _08958_ (.A1(\sha256cu.m_out_digest.e_in[10] ),
    .A2(_02070_),
    .B1(_03449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00233_));
 sky130_fd_sc_hd__or2b_1 _08959_ (.A(_03437_),
    .B_N(_03436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03450_));
 sky130_fd_sc_hd__nand2_1 _08960_ (.A(_03438_),
    .B(_03439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03451_));
 sky130_fd_sc_hd__nor2_1 _08961_ (.A(\sha256cu.m_out_digest.h_in[11] ),
    .B(\sha256cu.m_out_digest.d_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03452_));
 sky130_fd_sc_hd__and2_1 _08962_ (.A(\sha256cu.m_out_digest.h_in[11] ),
    .B(\sha256cu.m_out_digest.d_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03453_));
 sky130_fd_sc_hd__nor2_1 _08963_ (.A(_03452_),
    .B(_03453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03454_));
 sky130_fd_sc_hd__xnor2_1 _08964_ (.A(_02417_),
    .B(_03454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03455_));
 sky130_fd_sc_hd__a21boi_1 _08965_ (.A1(_02380_),
    .A2(_03423_),
    .B1_N(_03424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03456_));
 sky130_fd_sc_hd__xnor2_1 _08966_ (.A(_03455_),
    .B(_03456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03457_));
 sky130_fd_sc_hd__or2_1 _08967_ (.A(\sha256cu.iter_processing.w[11] ),
    .B(_02413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03458_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(\sha256cu.iter_processing.w[11] ),
    .B(_02413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03459_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_03458_),
    .B(_03459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03460_));
 sky130_fd_sc_hd__xor2_1 _08970_ (.A(\sha256cu.K[11] ),
    .B(_03460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03461_));
 sky130_fd_sc_hd__nor2_1 _08971_ (.A(_03457_),
    .B(_03461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03462_));
 sky130_fd_sc_hd__and2_1 _08972_ (.A(_03457_),
    .B(_03461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03463_));
 sky130_fd_sc_hd__nor2_1 _08973_ (.A(_03462_),
    .B(_03463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03464_));
 sky130_fd_sc_hd__o21ba_1 _08974_ (.A1(_03430_),
    .A2(_03435_),
    .B1_N(_03428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03465_));
 sky130_fd_sc_hd__xnor2_1 _08975_ (.A(_03464_),
    .B(_03465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03466_));
 sky130_fd_sc_hd__o21ai_1 _08976_ (.A1(_03431_),
    .A2(_03434_),
    .B1(_03433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03467_));
 sky130_fd_sc_hd__xnor2_1 _08977_ (.A(_03466_),
    .B(_03467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03468_));
 sky130_fd_sc_hd__and3_1 _08978_ (.A(_03450_),
    .B(_03451_),
    .C(_03468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03469_));
 sky130_fd_sc_hd__a21oi_1 _08979_ (.A1(_03450_),
    .A2(_03451_),
    .B1(_03468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03470_));
 sky130_fd_sc_hd__nor2_1 _08980_ (.A(_03469_),
    .B(_03470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03471_));
 sky130_fd_sc_hd__a21oi_1 _08981_ (.A1(_03441_),
    .A2(_03448_),
    .B1(_03471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03472_));
 sky130_fd_sc_hd__a31o_1 _08982_ (.A1(_03441_),
    .A2(_03448_),
    .A3(_03471_),
    .B1(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03473_));
 sky130_fd_sc_hd__or2_1 _08983_ (.A(\sha256cu.m_out_digest.e_in[11] ),
    .B(_02440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03474_));
 sky130_fd_sc_hd__o211a_1 _08984_ (.A1(_03472_),
    .A2(_03473_),
    .B1(_03474_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00234_));
 sky130_fd_sc_hd__nor2_1 _08985_ (.A(_03455_),
    .B(_03456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03475_));
 sky130_fd_sc_hd__nor2_1 _08986_ (.A(\sha256cu.m_out_digest.h_in[12] ),
    .B(\sha256cu.m_out_digest.d_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03476_));
 sky130_fd_sc_hd__and2_1 _08987_ (.A(\sha256cu.m_out_digest.h_in[12] ),
    .B(\sha256cu.m_out_digest.d_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03477_));
 sky130_fd_sc_hd__nor2_1 _08988_ (.A(_03476_),
    .B(_03477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03478_));
 sky130_fd_sc_hd__xnor2_1 _08989_ (.A(_02450_),
    .B(_03478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03479_));
 sky130_fd_sc_hd__a21oi_1 _08990_ (.A1(_02417_),
    .A2(_03454_),
    .B1(_03453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03480_));
 sky130_fd_sc_hd__xnor2_1 _08991_ (.A(_03479_),
    .B(_03480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03481_));
 sky130_fd_sc_hd__nor2_1 _08992_ (.A(\sha256cu.iter_processing.w[12] ),
    .B(_02446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03482_));
 sky130_fd_sc_hd__and2_1 _08993_ (.A(\sha256cu.iter_processing.w[12] ),
    .B(_02446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03483_));
 sky130_fd_sc_hd__nor2_1 _08994_ (.A(_03482_),
    .B(_03483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03484_));
 sky130_fd_sc_hd__xnor2_1 _08995_ (.A(\sha256cu.K[12] ),
    .B(_03484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03485_));
 sky130_fd_sc_hd__nor2_1 _08996_ (.A(_03481_),
    .B(_03485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03486_));
 sky130_fd_sc_hd__and2_1 _08997_ (.A(_03481_),
    .B(_03485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03487_));
 sky130_fd_sc_hd__nor2_1 _08998_ (.A(_03486_),
    .B(_03487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03488_));
 sky130_fd_sc_hd__o21ai_1 _08999_ (.A1(_03475_),
    .A2(_03462_),
    .B1(_03488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03489_));
 sky130_fd_sc_hd__or3_1 _09000_ (.A(_03475_),
    .B(_03462_),
    .C(_03488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03490_));
 sky130_fd_sc_hd__and2_1 _09001_ (.A(_03489_),
    .B(_03490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03491_));
 sky130_fd_sc_hd__a21bo_1 _09002_ (.A1(\sha256cu.K[11] ),
    .A2(_03458_),
    .B1_N(_03459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03492_));
 sky130_fd_sc_hd__xor2_1 _09003_ (.A(_03491_),
    .B(_03492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03493_));
 sky130_fd_sc_hd__or3_1 _09004_ (.A(_03462_),
    .B(_03463_),
    .C(_03465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03494_));
 sky130_fd_sc_hd__a21bo_1 _09005_ (.A1(_03466_),
    .A2(_03467_),
    .B1_N(_03494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03495_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(_03493_),
    .B(_03495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03496_));
 sky130_fd_sc_hd__or2_1 _09007_ (.A(_03493_),
    .B(_03495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03497_));
 sky130_fd_sc_hd__nand2_1 _09008_ (.A(_03496_),
    .B(_03497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03498_));
 sky130_fd_sc_hd__nand2_1 _09009_ (.A(_03443_),
    .B(_03471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03499_));
 sky130_fd_sc_hd__nor2_1 _09010_ (.A(_03441_),
    .B(_03469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03500_));
 sky130_fd_sc_hd__a311oi_1 _09011_ (.A1(_03443_),
    .A2(_03447_),
    .A3(_03471_),
    .B1(_03500_),
    .C1(_03470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03501_));
 sky130_fd_sc_hd__o31a_2 _09012_ (.A1(_03391_),
    .A2(_03444_),
    .A3(_03499_),
    .B1(_03501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03502_));
 sky130_fd_sc_hd__or2_1 _09013_ (.A(_03498_),
    .B(_03502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03503_));
 sky130_fd_sc_hd__a21oi_1 _09014_ (.A1(_03498_),
    .A2(_03502_),
    .B1(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03504_));
 sky130_fd_sc_hd__a221o_1 _09015_ (.A1(\sha256cu.m_out_digest.e_in[12] ),
    .A2(_02732_),
    .B1(_03503_),
    .B2(_03504_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00235_));
 sky130_fd_sc_hd__nand2_1 _09016_ (.A(_03491_),
    .B(_03492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03505_));
 sky130_fd_sc_hd__nor2_1 _09017_ (.A(_03479_),
    .B(_03480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03506_));
 sky130_fd_sc_hd__nor2_1 _09018_ (.A(\sha256cu.m_out_digest.h_in[13] ),
    .B(\sha256cu.m_out_digest.d_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03507_));
 sky130_fd_sc_hd__and2_1 _09019_ (.A(\sha256cu.m_out_digest.h_in[13] ),
    .B(\sha256cu.m_out_digest.d_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03508_));
 sky130_fd_sc_hd__nor2_1 _09020_ (.A(_03507_),
    .B(_03508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03509_));
 sky130_fd_sc_hd__xnor2_1 _09021_ (.A(_02492_),
    .B(_03509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03510_));
 sky130_fd_sc_hd__a21oi_1 _09022_ (.A1(_02450_),
    .A2(_03478_),
    .B1(_03477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03511_));
 sky130_fd_sc_hd__xnor2_1 _09023_ (.A(_03510_),
    .B(_03511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03512_));
 sky130_fd_sc_hd__nor2_1 _09024_ (.A(\sha256cu.iter_processing.w[13] ),
    .B(_02488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03513_));
 sky130_fd_sc_hd__and2_1 _09025_ (.A(\sha256cu.iter_processing.w[13] ),
    .B(_02488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03514_));
 sky130_fd_sc_hd__nor2_1 _09026_ (.A(_03513_),
    .B(_03514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03515_));
 sky130_fd_sc_hd__xnor2_1 _09027_ (.A(\sha256cu.K[13] ),
    .B(_03515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03516_));
 sky130_fd_sc_hd__nor2_1 _09028_ (.A(_03512_),
    .B(_03516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03517_));
 sky130_fd_sc_hd__and2_1 _09029_ (.A(_03512_),
    .B(_03516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03518_));
 sky130_fd_sc_hd__nor2_1 _09030_ (.A(_03517_),
    .B(_03518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03519_));
 sky130_fd_sc_hd__o21ai_1 _09031_ (.A1(_03506_),
    .A2(_03486_),
    .B1(_03519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03520_));
 sky130_fd_sc_hd__or3_1 _09032_ (.A(_03506_),
    .B(_03486_),
    .C(_03519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03521_));
 sky130_fd_sc_hd__and2_1 _09033_ (.A(_03520_),
    .B(_03521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03522_));
 sky130_fd_sc_hd__a21o_1 _09034_ (.A1(\sha256cu.K[12] ),
    .A2(_03484_),
    .B1(_03483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03523_));
 sky130_fd_sc_hd__xnor2_1 _09035_ (.A(_03522_),
    .B(_03523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03524_));
 sky130_fd_sc_hd__and3_1 _09036_ (.A(_03489_),
    .B(_03505_),
    .C(_03524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03525_));
 sky130_fd_sc_hd__a21o_1 _09037_ (.A1(_03489_),
    .A2(_03505_),
    .B1(_03524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03526_));
 sky130_fd_sc_hd__and2b_1 _09038_ (.A_N(_03525_),
    .B(_03526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03527_));
 sky130_fd_sc_hd__a21oi_1 _09039_ (.A1(_03496_),
    .A2(_03503_),
    .B1(_03527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03528_));
 sky130_fd_sc_hd__a31o_1 _09040_ (.A1(_03496_),
    .A2(_03503_),
    .A3(_03527_),
    .B1(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03529_));
 sky130_fd_sc_hd__or2_1 _09041_ (.A(\sha256cu.m_out_digest.e_in[13] ),
    .B(_02440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03530_));
 sky130_fd_sc_hd__o211a_1 _09042_ (.A1(_03528_),
    .A2(_03529_),
    .B1(_03530_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00236_));
 sky130_fd_sc_hd__nand2_1 _09043_ (.A(_03522_),
    .B(_03523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03531_));
 sky130_fd_sc_hd__nor2_1 _09044_ (.A(_03510_),
    .B(_03511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03532_));
 sky130_fd_sc_hd__or2_1 _09045_ (.A(\sha256cu.m_out_digest.h_in[14] ),
    .B(\sha256cu.m_out_digest.d_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03533_));
 sky130_fd_sc_hd__nand2_1 _09046_ (.A(\sha256cu.m_out_digest.h_in[14] ),
    .B(\sha256cu.m_out_digest.d_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03534_));
 sky130_fd_sc_hd__nand2_1 _09047_ (.A(_03533_),
    .B(_03534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03535_));
 sky130_fd_sc_hd__xor2_1 _09048_ (.A(_02525_),
    .B(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03536_));
 sky130_fd_sc_hd__a21oi_1 _09049_ (.A1(_02492_),
    .A2(_03509_),
    .B1(_03508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03537_));
 sky130_fd_sc_hd__or2_1 _09050_ (.A(_03536_),
    .B(_03537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03538_));
 sky130_fd_sc_hd__nand2_1 _09051_ (.A(_03536_),
    .B(_03537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03539_));
 sky130_fd_sc_hd__nand2_1 _09052_ (.A(_03538_),
    .B(_03539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03540_));
 sky130_fd_sc_hd__nor2_1 _09053_ (.A(\sha256cu.iter_processing.w[14] ),
    .B(_02521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03541_));
 sky130_fd_sc_hd__and2_1 _09054_ (.A(\sha256cu.iter_processing.w[14] ),
    .B(_02521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03542_));
 sky130_fd_sc_hd__nor2_1 _09055_ (.A(_03541_),
    .B(_03542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03543_));
 sky130_fd_sc_hd__xnor2_1 _09056_ (.A(\sha256cu.K[14] ),
    .B(_03543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03544_));
 sky130_fd_sc_hd__xor2_1 _09057_ (.A(_03540_),
    .B(_03544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03545_));
 sky130_fd_sc_hd__o21ai_1 _09058_ (.A1(_03532_),
    .A2(_03517_),
    .B1(_03545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03546_));
 sky130_fd_sc_hd__or3_1 _09059_ (.A(_03532_),
    .B(_03517_),
    .C(_03545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03547_));
 sky130_fd_sc_hd__and2_1 _09060_ (.A(_03546_),
    .B(_03547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03548_));
 sky130_fd_sc_hd__a21o_1 _09061_ (.A1(\sha256cu.K[13] ),
    .A2(_03515_),
    .B1(_03514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03549_));
 sky130_fd_sc_hd__xnor2_1 _09062_ (.A(_03548_),
    .B(_03549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03550_));
 sky130_fd_sc_hd__a21o_1 _09063_ (.A1(_03520_),
    .A2(_03531_),
    .B1(_03550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03551_));
 sky130_fd_sc_hd__nand3_1 _09064_ (.A(_03520_),
    .B(_03531_),
    .C(_03550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03552_));
 sky130_fd_sc_hd__and2_1 _09065_ (.A(_03551_),
    .B(_03552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03553_));
 sky130_fd_sc_hd__or2b_1 _09066_ (.A(_03498_),
    .B_N(_03527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03554_));
 sky130_fd_sc_hd__a21oi_1 _09067_ (.A1(_03496_),
    .A2(_03526_),
    .B1(_03525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03555_));
 sky130_fd_sc_hd__o21bai_1 _09068_ (.A1(_03502_),
    .A2(_03554_),
    .B1_N(_03555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03556_));
 sky130_fd_sc_hd__nand2_1 _09069_ (.A(_03553_),
    .B(_03556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03557_));
 sky130_fd_sc_hd__o21a_1 _09070_ (.A1(_03553_),
    .A2(_03556_),
    .B1(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03558_));
 sky130_fd_sc_hd__a221o_1 _09071_ (.A1(\sha256cu.m_out_digest.e_in[14] ),
    .A2(_02732_),
    .B1(_03557_),
    .B2(_03558_),
    .C1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00237_));
 sky130_fd_sc_hd__clkbuf_4 _09072_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03559_));
 sky130_fd_sc_hd__nand2_1 _09073_ (.A(_03548_),
    .B(_03549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03560_));
 sky130_fd_sc_hd__or2_1 _09074_ (.A(\sha256cu.m_out_digest.h_in[15] ),
    .B(\sha256cu.m_out_digest.d_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_1 _09075_ (.A(\sha256cu.m_out_digest.h_in[15] ),
    .B(\sha256cu.m_out_digest.d_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03562_));
 sky130_fd_sc_hd__nand2_1 _09076_ (.A(_03561_),
    .B(_03562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03563_));
 sky130_fd_sc_hd__xor2_1 _09077_ (.A(_02565_),
    .B(_03563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03564_));
 sky130_fd_sc_hd__o21a_1 _09078_ (.A1(_02526_),
    .A2(_03535_),
    .B1(_03534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03565_));
 sky130_fd_sc_hd__nor2_1 _09079_ (.A(_03564_),
    .B(_03565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03566_));
 sky130_fd_sc_hd__and2_1 _09080_ (.A(_03564_),
    .B(_03565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03567_));
 sky130_fd_sc_hd__or2_1 _09081_ (.A(_03566_),
    .B(_03567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03568_));
 sky130_fd_sc_hd__or2_1 _09082_ (.A(\sha256cu.iter_processing.w[15] ),
    .B(_02561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03569_));
 sky130_fd_sc_hd__and2_1 _09083_ (.A(\sha256cu.iter_processing.w[15] ),
    .B(_02561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03570_));
 sky130_fd_sc_hd__inv_2 _09084_ (.A(_03570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03571_));
 sky130_fd_sc_hd__nand2_1 _09085_ (.A(_03569_),
    .B(_03571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03572_));
 sky130_fd_sc_hd__xor2_1 _09086_ (.A(\sha256cu.K[15] ),
    .B(_03572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03573_));
 sky130_fd_sc_hd__xor2_1 _09087_ (.A(_03568_),
    .B(_03573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03574_));
 sky130_fd_sc_hd__o21a_1 _09088_ (.A1(_03540_),
    .A2(_03544_),
    .B1(_03538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03575_));
 sky130_fd_sc_hd__xnor2_1 _09089_ (.A(_03574_),
    .B(_03575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03576_));
 sky130_fd_sc_hd__a21o_1 _09090_ (.A1(\sha256cu.K[14] ),
    .A2(_03543_),
    .B1(_03542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03577_));
 sky130_fd_sc_hd__xnor2_1 _09091_ (.A(_03576_),
    .B(_03577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03578_));
 sky130_fd_sc_hd__and3_1 _09092_ (.A(_03546_),
    .B(_03560_),
    .C(_03578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03579_));
 sky130_fd_sc_hd__a21oi_1 _09093_ (.A1(_03546_),
    .A2(_03560_),
    .B1(_03578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03580_));
 sky130_fd_sc_hd__nor2_1 _09094_ (.A(_03579_),
    .B(_03580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03581_));
 sky130_fd_sc_hd__and3_1 _09095_ (.A(_03551_),
    .B(_03557_),
    .C(_03581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03582_));
 sky130_fd_sc_hd__a21oi_1 _09096_ (.A1(_03551_),
    .A2(_03557_),
    .B1(_03581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03583_));
 sky130_fd_sc_hd__or2_1 _09097_ (.A(_03582_),
    .B(_03583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03584_));
 sky130_fd_sc_hd__a22o_1 _09098_ (.A1(\sha256cu.m_out_digest.e_in[15] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(_03584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00238_));
 sky130_fd_sc_hd__or2_1 _09099_ (.A(\sha256cu.m_out_digest.h_in[16] ),
    .B(\sha256cu.m_out_digest.d_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03585_));
 sky130_fd_sc_hd__nand2_1 _09100_ (.A(\sha256cu.m_out_digest.h_in[16] ),
    .B(\sha256cu.m_out_digest.d_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(_03585_),
    .B(_03586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03587_));
 sky130_fd_sc_hd__xor2_1 _09102_ (.A(_02599_),
    .B(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03588_));
 sky130_fd_sc_hd__a21boi_1 _09103_ (.A1(_02565_),
    .A2(_03561_),
    .B1_N(_03562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03589_));
 sky130_fd_sc_hd__nor2_1 _09104_ (.A(_03588_),
    .B(_03589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03590_));
 sky130_fd_sc_hd__and2_1 _09105_ (.A(_03588_),
    .B(_03589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03591_));
 sky130_fd_sc_hd__or2_1 _09106_ (.A(_03590_),
    .B(_03591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03592_));
 sky130_fd_sc_hd__nor2_1 _09107_ (.A(\sha256cu.iter_processing.w[16] ),
    .B(_02595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03593_));
 sky130_fd_sc_hd__and2_1 _09108_ (.A(\sha256cu.iter_processing.w[16] ),
    .B(_02595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03594_));
 sky130_fd_sc_hd__nor2_1 _09109_ (.A(_03593_),
    .B(_03594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03595_));
 sky130_fd_sc_hd__xnor2_1 _09110_ (.A(\sha256cu.K[16] ),
    .B(_03595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03596_));
 sky130_fd_sc_hd__nor2_1 _09111_ (.A(_03592_),
    .B(_03596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03597_));
 sky130_fd_sc_hd__and2_1 _09112_ (.A(_03592_),
    .B(_03596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03598_));
 sky130_fd_sc_hd__nor2_1 _09113_ (.A(_03597_),
    .B(_03598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03599_));
 sky130_fd_sc_hd__o21ba_1 _09114_ (.A1(_03567_),
    .A2(_03573_),
    .B1_N(_03566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03600_));
 sky130_fd_sc_hd__xnor2_1 _09115_ (.A(_03599_),
    .B(_03600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03601_));
 sky130_fd_sc_hd__a21o_1 _09116_ (.A1(\sha256cu.K[15] ),
    .A2(_03569_),
    .B1(_03570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03602_));
 sky130_fd_sc_hd__xor2_1 _09117_ (.A(_03601_),
    .B(_03602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03603_));
 sky130_fd_sc_hd__or2b_1 _09118_ (.A(_03575_),
    .B_N(_03574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03604_));
 sky130_fd_sc_hd__a21bo_1 _09119_ (.A1(_03576_),
    .A2(_03577_),
    .B1_N(_03604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03605_));
 sky130_fd_sc_hd__nand2_1 _09120_ (.A(_03603_),
    .B(_03605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03606_));
 sky130_fd_sc_hd__or2_1 _09121_ (.A(_03603_),
    .B(_03605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03607_));
 sky130_fd_sc_hd__and2_1 _09122_ (.A(_03606_),
    .B(_03607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03608_));
 sky130_fd_sc_hd__nand2_1 _09123_ (.A(_03553_),
    .B(_03581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03609_));
 sky130_fd_sc_hd__nor2_1 _09124_ (.A(_03551_),
    .B(_03579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03610_));
 sky130_fd_sc_hd__a311oi_1 _09125_ (.A1(_03553_),
    .A2(_03555_),
    .A3(_03581_),
    .B1(_03610_),
    .C1(_03580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03611_));
 sky130_fd_sc_hd__o31a_1 _09126_ (.A1(_03502_),
    .A2(_03554_),
    .A3(_03609_),
    .B1(_03611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03612_));
 sky130_fd_sc_hd__xnor2_1 _09127_ (.A(_03608_),
    .B(_03612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03613_));
 sky130_fd_sc_hd__or2_1 _09128_ (.A(\sha256cu.m_out_digest.e_in[16] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03614_));
 sky130_fd_sc_hd__o211a_1 _09129_ (.A1(_02040_),
    .A2(_03613_),
    .B1(_03614_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00239_));
 sky130_fd_sc_hd__or3_1 _09130_ (.A(_03597_),
    .B(_03598_),
    .C(_03600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03615_));
 sky130_fd_sc_hd__nand2_1 _09131_ (.A(_03601_),
    .B(_03602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03616_));
 sky130_fd_sc_hd__or2_1 _09132_ (.A(\sha256cu.m_out_digest.h_in[17] ),
    .B(\sha256cu.m_out_digest.d_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03617_));
 sky130_fd_sc_hd__nand2_1 _09133_ (.A(\sha256cu.m_out_digest.h_in[17] ),
    .B(\sha256cu.m_out_digest.d_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _09134_ (.A(_03617_),
    .B(_03618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03619_));
 sky130_fd_sc_hd__xor2_1 _09135_ (.A(_02643_),
    .B(_03619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03620_));
 sky130_fd_sc_hd__a21boi_1 _09136_ (.A1(_02599_),
    .A2(_03585_),
    .B1_N(_03586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03621_));
 sky130_fd_sc_hd__xnor2_1 _09137_ (.A(_03620_),
    .B(_03621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03622_));
 sky130_fd_sc_hd__nor2_1 _09138_ (.A(\sha256cu.iter_processing.w[17] ),
    .B(_02639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03623_));
 sky130_fd_sc_hd__and2_1 _09139_ (.A(\sha256cu.iter_processing.w[17] ),
    .B(_02639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03624_));
 sky130_fd_sc_hd__nor2_1 _09140_ (.A(_03623_),
    .B(_03624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03625_));
 sky130_fd_sc_hd__xnor2_1 _09141_ (.A(\sha256cu.K[17] ),
    .B(_03625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03626_));
 sky130_fd_sc_hd__nor2_1 _09142_ (.A(_03622_),
    .B(_03626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03627_));
 sky130_fd_sc_hd__and2_1 _09143_ (.A(_03622_),
    .B(_03626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03628_));
 sky130_fd_sc_hd__nor2_1 _09144_ (.A(_03627_),
    .B(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03629_));
 sky130_fd_sc_hd__o21ai_1 _09145_ (.A1(_03590_),
    .A2(_03597_),
    .B1(_03629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03630_));
 sky130_fd_sc_hd__or3_1 _09146_ (.A(_03590_),
    .B(_03597_),
    .C(_03629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03631_));
 sky130_fd_sc_hd__and2_1 _09147_ (.A(_03630_),
    .B(_03631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03632_));
 sky130_fd_sc_hd__a21o_1 _09148_ (.A1(\sha256cu.K[16] ),
    .A2(_03595_),
    .B1(_03594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03633_));
 sky130_fd_sc_hd__xnor2_1 _09149_ (.A(_03632_),
    .B(_03633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03634_));
 sky130_fd_sc_hd__and3_1 _09150_ (.A(_03615_),
    .B(_03616_),
    .C(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03635_));
 sky130_fd_sc_hd__a21o_1 _09151_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03636_));
 sky130_fd_sc_hd__and2b_1 _09152_ (.A_N(_03635_),
    .B(_03636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03637_));
 sky130_fd_sc_hd__inv_2 _09153_ (.A(_03612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03638_));
 sky130_fd_sc_hd__a21bo_1 _09154_ (.A1(_03608_),
    .A2(_03638_),
    .B1_N(_03606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03639_));
 sky130_fd_sc_hd__xnor2_1 _09155_ (.A(_03637_),
    .B(_03639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03640_));
 sky130_fd_sc_hd__nor2_1 _09156_ (.A(_02069_),
    .B(_03640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03641_));
 sky130_fd_sc_hd__a211o_1 _09157_ (.A1(\sha256cu.m_out_digest.e_in[17] ),
    .A2(_02040_),
    .B1(_03641_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00240_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(_03632_),
    .B(_03633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03642_));
 sky130_fd_sc_hd__nor2_1 _09159_ (.A(_03620_),
    .B(_03621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03643_));
 sky130_fd_sc_hd__or2_1 _09160_ (.A(\sha256cu.m_out_digest.h_in[18] ),
    .B(\sha256cu.m_out_digest.d_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03644_));
 sky130_fd_sc_hd__nand2_1 _09161_ (.A(\sha256cu.m_out_digest.h_in[18] ),
    .B(\sha256cu.m_out_digest.d_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03645_));
 sky130_fd_sc_hd__nand2_1 _09162_ (.A(_03644_),
    .B(_03645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03646_));
 sky130_fd_sc_hd__xor2_1 _09163_ (.A(_02675_),
    .B(_03646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03647_));
 sky130_fd_sc_hd__a21boi_1 _09164_ (.A1(_02643_),
    .A2(_03617_),
    .B1_N(_03618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03648_));
 sky130_fd_sc_hd__xnor2_1 _09165_ (.A(_03647_),
    .B(_03648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03649_));
 sky130_fd_sc_hd__nor2_1 _09166_ (.A(\sha256cu.iter_processing.w[18] ),
    .B(_02671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03650_));
 sky130_fd_sc_hd__and2_1 _09167_ (.A(\sha256cu.iter_processing.w[18] ),
    .B(_02671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03651_));
 sky130_fd_sc_hd__nor2_1 _09168_ (.A(_03650_),
    .B(_03651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03652_));
 sky130_fd_sc_hd__xnor2_1 _09169_ (.A(\sha256cu.K[18] ),
    .B(_03652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03653_));
 sky130_fd_sc_hd__nor2_1 _09170_ (.A(_03649_),
    .B(_03653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03654_));
 sky130_fd_sc_hd__and2_1 _09171_ (.A(_03649_),
    .B(_03653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03655_));
 sky130_fd_sc_hd__nor2_1 _09172_ (.A(_03654_),
    .B(_03655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03656_));
 sky130_fd_sc_hd__o21ai_1 _09173_ (.A1(_03643_),
    .A2(_03627_),
    .B1(_03656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03657_));
 sky130_fd_sc_hd__or3_1 _09174_ (.A(_03643_),
    .B(_03627_),
    .C(_03656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03658_));
 sky130_fd_sc_hd__and2_1 _09175_ (.A(_03657_),
    .B(_03658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03659_));
 sky130_fd_sc_hd__a21o_1 _09176_ (.A1(\sha256cu.K[17] ),
    .A2(_03625_),
    .B1(_03624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03660_));
 sky130_fd_sc_hd__xnor2_1 _09177_ (.A(_03659_),
    .B(_03660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03661_));
 sky130_fd_sc_hd__a21oi_1 _09178_ (.A1(_03630_),
    .A2(_03642_),
    .B1(_03661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03662_));
 sky130_fd_sc_hd__and3_1 _09179_ (.A(_03630_),
    .B(_03642_),
    .C(_03661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03663_));
 sky130_fd_sc_hd__nor2_1 _09180_ (.A(_03662_),
    .B(_03663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03664_));
 sky130_fd_sc_hd__a21oi_1 _09181_ (.A1(_03606_),
    .A2(_03636_),
    .B1(_03635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03665_));
 sky130_fd_sc_hd__a31o_1 _09182_ (.A1(_03608_),
    .A2(_03638_),
    .A3(_03637_),
    .B1(_03665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03666_));
 sky130_fd_sc_hd__xnor2_1 _09183_ (.A(_03664_),
    .B(_03666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03667_));
 sky130_fd_sc_hd__nor2_1 _09184_ (.A(_02069_),
    .B(_03667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03668_));
 sky130_fd_sc_hd__a211o_1 _09185_ (.A1(\sha256cu.m_out_digest.e_in[18] ),
    .A2(_02040_),
    .B1(_03668_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00241_));
 sky130_fd_sc_hd__nand2_1 _09186_ (.A(_03659_),
    .B(_03660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03669_));
 sky130_fd_sc_hd__nor2_1 _09187_ (.A(_03647_),
    .B(_03648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03670_));
 sky130_fd_sc_hd__or2_1 _09188_ (.A(\sha256cu.m_out_digest.h_in[19] ),
    .B(\sha256cu.m_out_digest.d_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03671_));
 sky130_fd_sc_hd__nand2_1 _09189_ (.A(\sha256cu.m_out_digest.h_in[19] ),
    .B(\sha256cu.m_out_digest.d_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_1 _09190_ (.A(_03671_),
    .B(_03672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03673_));
 sky130_fd_sc_hd__xor2_1 _09191_ (.A(_02712_),
    .B(_03673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03674_));
 sky130_fd_sc_hd__a21boi_1 _09192_ (.A1(_02675_),
    .A2(_03644_),
    .B1_N(_03645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03675_));
 sky130_fd_sc_hd__xnor2_1 _09193_ (.A(_03674_),
    .B(_03675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03676_));
 sky130_fd_sc_hd__or2_1 _09194_ (.A(\sha256cu.iter_processing.w[19] ),
    .B(_02708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03677_));
 sky130_fd_sc_hd__nand2_1 _09195_ (.A(\sha256cu.iter_processing.w[19] ),
    .B(_02708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03678_));
 sky130_fd_sc_hd__nand2_1 _09196_ (.A(_03677_),
    .B(_03678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03679_));
 sky130_fd_sc_hd__xor2_1 _09197_ (.A(\sha256cu.K[19] ),
    .B(_03679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03680_));
 sky130_fd_sc_hd__nor2_1 _09198_ (.A(_03676_),
    .B(_03680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03681_));
 sky130_fd_sc_hd__and2_1 _09199_ (.A(_03676_),
    .B(_03680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03682_));
 sky130_fd_sc_hd__nor2_1 _09200_ (.A(_03681_),
    .B(_03682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03683_));
 sky130_fd_sc_hd__o21a_1 _09201_ (.A1(_03670_),
    .A2(_03654_),
    .B1(_03683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03684_));
 sky130_fd_sc_hd__nor3_1 _09202_ (.A(_03670_),
    .B(_03654_),
    .C(_03683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03685_));
 sky130_fd_sc_hd__nor2_1 _09203_ (.A(_03684_),
    .B(_03685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03686_));
 sky130_fd_sc_hd__a21o_1 _09204_ (.A1(\sha256cu.K[18] ),
    .A2(_03652_),
    .B1(_03651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03687_));
 sky130_fd_sc_hd__xnor2_1 _09205_ (.A(_03686_),
    .B(_03687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03688_));
 sky130_fd_sc_hd__and3_1 _09206_ (.A(_03657_),
    .B(_03669_),
    .C(_03688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03689_));
 sky130_fd_sc_hd__a21oi_1 _09207_ (.A1(_03657_),
    .A2(_03669_),
    .B1(_03688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03690_));
 sky130_fd_sc_hd__nor2_1 _09208_ (.A(_03689_),
    .B(_03690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03691_));
 sky130_fd_sc_hd__a21o_1 _09209_ (.A1(_03664_),
    .A2(_03666_),
    .B1(_03662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03692_));
 sky130_fd_sc_hd__nor2_1 _09210_ (.A(_03691_),
    .B(_03692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03693_));
 sky130_fd_sc_hd__a211oi_1 _09211_ (.A1(_03691_),
    .A2(_03692_),
    .B1(_03693_),
    .C1(_02732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03694_));
 sky130_fd_sc_hd__a211o_1 _09212_ (.A1(\sha256cu.m_out_digest.e_in[19] ),
    .A2(_02040_),
    .B1(_03694_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00242_));
 sky130_fd_sc_hd__nor2_1 _09213_ (.A(_03674_),
    .B(_03675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03695_));
 sky130_fd_sc_hd__or2_1 _09214_ (.A(\sha256cu.m_out_digest.h_in[20] ),
    .B(\sha256cu.m_out_digest.d_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03696_));
 sky130_fd_sc_hd__nand2_1 _09215_ (.A(\sha256cu.m_out_digest.h_in[20] ),
    .B(\sha256cu.m_out_digest.d_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03697_));
 sky130_fd_sc_hd__nand2_1 _09216_ (.A(_03696_),
    .B(_03697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03698_));
 sky130_fd_sc_hd__xor2_1 _09217_ (.A(_02747_),
    .B(_03698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03699_));
 sky130_fd_sc_hd__a21boi_1 _09218_ (.A1(_02712_),
    .A2(_03671_),
    .B1_N(_03672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03700_));
 sky130_fd_sc_hd__nor2_1 _09219_ (.A(_03699_),
    .B(_03700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03701_));
 sky130_fd_sc_hd__and2_1 _09220_ (.A(_03699_),
    .B(_03700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03702_));
 sky130_fd_sc_hd__or2_1 _09221_ (.A(_03701_),
    .B(_03702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03703_));
 sky130_fd_sc_hd__nor2_1 _09222_ (.A(\sha256cu.iter_processing.w[20] ),
    .B(_02740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03704_));
 sky130_fd_sc_hd__and2_1 _09223_ (.A(\sha256cu.iter_processing.w[20] ),
    .B(_02740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03705_));
 sky130_fd_sc_hd__nor2_1 _09224_ (.A(_03704_),
    .B(_03705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03706_));
 sky130_fd_sc_hd__xnor2_1 _09225_ (.A(\sha256cu.K[20] ),
    .B(_03706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03707_));
 sky130_fd_sc_hd__nor2_1 _09226_ (.A(_03703_),
    .B(_03707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03708_));
 sky130_fd_sc_hd__and2_1 _09227_ (.A(_03703_),
    .B(_03707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03709_));
 sky130_fd_sc_hd__nor2_1 _09228_ (.A(_03708_),
    .B(_03709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03710_));
 sky130_fd_sc_hd__o21ai_1 _09229_ (.A1(_03695_),
    .A2(_03681_),
    .B1(_03710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03711_));
 sky130_fd_sc_hd__or3_1 _09230_ (.A(_03695_),
    .B(_03681_),
    .C(_03710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03712_));
 sky130_fd_sc_hd__and2_1 _09231_ (.A(_03711_),
    .B(_03712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03713_));
 sky130_fd_sc_hd__a21bo_1 _09232_ (.A1(\sha256cu.K[19] ),
    .A2(_03677_),
    .B1_N(_03678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03714_));
 sky130_fd_sc_hd__xor2_1 _09233_ (.A(_03713_),
    .B(_03714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03715_));
 sky130_fd_sc_hd__a21o_1 _09234_ (.A1(_03686_),
    .A2(_03687_),
    .B1(_03684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03716_));
 sky130_fd_sc_hd__nand2_1 _09235_ (.A(_03715_),
    .B(_03716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03717_));
 sky130_fd_sc_hd__or2_1 _09236_ (.A(_03715_),
    .B(_03716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03718_));
 sky130_fd_sc_hd__and2_1 _09237_ (.A(_03717_),
    .B(_03718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03719_));
 sky130_fd_sc_hd__nand2_1 _09238_ (.A(_03608_),
    .B(_03637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03720_));
 sky130_fd_sc_hd__nand2_1 _09239_ (.A(_03664_),
    .B(_03691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03721_));
 sky130_fd_sc_hd__inv_2 _09240_ (.A(_03689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03722_));
 sky130_fd_sc_hd__a32o_1 _09241_ (.A1(_03664_),
    .A2(_03665_),
    .A3(_03691_),
    .B1(_03722_),
    .B2(_03662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03723_));
 sky130_fd_sc_hd__nor2_1 _09242_ (.A(_03690_),
    .B(_03723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03724_));
 sky130_fd_sc_hd__o31a_2 _09243_ (.A1(_03612_),
    .A2(_03720_),
    .A3(_03721_),
    .B1(_03724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03725_));
 sky130_fd_sc_hd__xnor2_1 _09244_ (.A(_03719_),
    .B(_03725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03726_));
 sky130_fd_sc_hd__or2_1 _09245_ (.A(\sha256cu.m_out_digest.e_in[20] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03727_));
 sky130_fd_sc_hd__o211a_1 _09246_ (.A1(_02040_),
    .A2(_03726_),
    .B1(_03727_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00243_));
 sky130_fd_sc_hd__nand2_1 _09247_ (.A(_03713_),
    .B(_03714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03728_));
 sky130_fd_sc_hd__or2_1 _09248_ (.A(\sha256cu.m_out_digest.h_in[21] ),
    .B(\sha256cu.m_out_digest.d_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03729_));
 sky130_fd_sc_hd__nand2_1 _09249_ (.A(\sha256cu.m_out_digest.h_in[21] ),
    .B(\sha256cu.m_out_digest.d_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03730_));
 sky130_fd_sc_hd__nand2_1 _09250_ (.A(_03729_),
    .B(_03730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03731_));
 sky130_fd_sc_hd__xor2_1 _09251_ (.A(_02777_),
    .B(_03731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03732_));
 sky130_fd_sc_hd__a21boi_1 _09252_ (.A1(_02747_),
    .A2(_03696_),
    .B1_N(_03697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03733_));
 sky130_fd_sc_hd__nor2_1 _09253_ (.A(_03732_),
    .B(_03733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03734_));
 sky130_fd_sc_hd__and2_1 _09254_ (.A(_03732_),
    .B(_03733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03735_));
 sky130_fd_sc_hd__or2_1 _09255_ (.A(_03734_),
    .B(_03735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03736_));
 sky130_fd_sc_hd__nor2_1 _09256_ (.A(\sha256cu.iter_processing.w[21] ),
    .B(_02785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03737_));
 sky130_fd_sc_hd__and2_1 _09257_ (.A(\sha256cu.iter_processing.w[21] ),
    .B(_02785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03738_));
 sky130_fd_sc_hd__nor2_1 _09258_ (.A(_03737_),
    .B(_03738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03739_));
 sky130_fd_sc_hd__xnor2_1 _09259_ (.A(\sha256cu.K[21] ),
    .B(_03739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03740_));
 sky130_fd_sc_hd__nor2_1 _09260_ (.A(_03736_),
    .B(_03740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03741_));
 sky130_fd_sc_hd__and2_1 _09261_ (.A(_03736_),
    .B(_03740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03742_));
 sky130_fd_sc_hd__nor2_1 _09262_ (.A(_03741_),
    .B(_03742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03743_));
 sky130_fd_sc_hd__o21ai_1 _09263_ (.A1(_03701_),
    .A2(_03708_),
    .B1(_03743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03744_));
 sky130_fd_sc_hd__or3_1 _09264_ (.A(_03701_),
    .B(_03708_),
    .C(_03743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03745_));
 sky130_fd_sc_hd__and2_1 _09265_ (.A(_03744_),
    .B(_03745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03746_));
 sky130_fd_sc_hd__a21o_1 _09266_ (.A1(\sha256cu.K[20] ),
    .A2(_03706_),
    .B1(_03705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03747_));
 sky130_fd_sc_hd__xnor2_1 _09267_ (.A(_03746_),
    .B(_03747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03748_));
 sky130_fd_sc_hd__and3_1 _09268_ (.A(_03711_),
    .B(_03728_),
    .C(_03748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03749_));
 sky130_fd_sc_hd__a21o_1 _09269_ (.A1(_03711_),
    .A2(_03728_),
    .B1(_03748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03750_));
 sky130_fd_sc_hd__and2b_1 _09270_ (.A_N(_03749_),
    .B(_03750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03751_));
 sky130_fd_sc_hd__inv_2 _09271_ (.A(_03725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03752_));
 sky130_fd_sc_hd__a21bo_1 _09272_ (.A1(_03719_),
    .A2(_03752_),
    .B1_N(_03717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03753_));
 sky130_fd_sc_hd__xor2_1 _09273_ (.A(_03751_),
    .B(_03753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03754_));
 sky130_fd_sc_hd__or2_1 _09274_ (.A(\sha256cu.m_out_digest.e_in[21] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03755_));
 sky130_fd_sc_hd__o211a_1 _09275_ (.A1(_02332_),
    .A2(_03754_),
    .B1(_03755_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00244_));
 sky130_fd_sc_hd__nand2_1 _09276_ (.A(_03746_),
    .B(_03747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03756_));
 sky130_fd_sc_hd__or2_1 _09277_ (.A(\sha256cu.m_out_digest.h_in[22] ),
    .B(\sha256cu.m_out_digest.d_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03757_));
 sky130_fd_sc_hd__nand2_1 _09278_ (.A(\sha256cu.m_out_digest.h_in[22] ),
    .B(\sha256cu.m_out_digest.d_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_1 _09279_ (.A(_03757_),
    .B(_03758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03759_));
 sky130_fd_sc_hd__xor2_1 _09280_ (.A(_02811_),
    .B(_03759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03760_));
 sky130_fd_sc_hd__a21boi_1 _09281_ (.A1(_02777_),
    .A2(_03729_),
    .B1_N(_03730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03761_));
 sky130_fd_sc_hd__nor2_1 _09282_ (.A(_03760_),
    .B(_03761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03762_));
 sky130_fd_sc_hd__and2_1 _09283_ (.A(_03760_),
    .B(_03761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03763_));
 sky130_fd_sc_hd__or2_1 _09284_ (.A(_03762_),
    .B(_03763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03764_));
 sky130_fd_sc_hd__nor2_1 _09285_ (.A(\sha256cu.iter_processing.w[22] ),
    .B(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03765_));
 sky130_fd_sc_hd__and2_1 _09286_ (.A(\sha256cu.iter_processing.w[22] ),
    .B(_02819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03766_));
 sky130_fd_sc_hd__nor2_1 _09287_ (.A(_03765_),
    .B(_03766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03767_));
 sky130_fd_sc_hd__xnor2_1 _09288_ (.A(\sha256cu.K[22] ),
    .B(_03767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03768_));
 sky130_fd_sc_hd__nor2_1 _09289_ (.A(_03764_),
    .B(_03768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03769_));
 sky130_fd_sc_hd__and2_1 _09290_ (.A(_03764_),
    .B(_03768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03770_));
 sky130_fd_sc_hd__nor2_1 _09291_ (.A(_03769_),
    .B(_03770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03771_));
 sky130_fd_sc_hd__o21ai_1 _09292_ (.A1(_03734_),
    .A2(_03741_),
    .B1(_03771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03772_));
 sky130_fd_sc_hd__or3_1 _09293_ (.A(_03734_),
    .B(_03741_),
    .C(_03771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03773_));
 sky130_fd_sc_hd__and2_1 _09294_ (.A(_03772_),
    .B(_03773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03774_));
 sky130_fd_sc_hd__a21o_1 _09295_ (.A1(\sha256cu.K[21] ),
    .A2(_03739_),
    .B1(_03738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03775_));
 sky130_fd_sc_hd__xnor2_1 _09296_ (.A(_03774_),
    .B(_03775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03776_));
 sky130_fd_sc_hd__a21o_1 _09297_ (.A1(_03744_),
    .A2(_03756_),
    .B1(_03776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03777_));
 sky130_fd_sc_hd__nand3_1 _09298_ (.A(_03744_),
    .B(_03756_),
    .C(_03776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03778_));
 sky130_fd_sc_hd__and2_1 _09299_ (.A(_03777_),
    .B(_03778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03779_));
 sky130_fd_sc_hd__nand2_1 _09300_ (.A(_03719_),
    .B(_03751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03780_));
 sky130_fd_sc_hd__nor2_1 _09301_ (.A(_03725_),
    .B(_03780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03781_));
 sky130_fd_sc_hd__a21oi_2 _09302_ (.A1(_03717_),
    .A2(_03750_),
    .B1(_03749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03782_));
 sky130_fd_sc_hd__or3_1 _09303_ (.A(_03779_),
    .B(_03781_),
    .C(_03782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03783_));
 sky130_fd_sc_hd__o21ai_1 _09304_ (.A1(_03781_),
    .A2(_03782_),
    .B1(_03779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03784_));
 sky130_fd_sc_hd__a32o_1 _09305_ (.A1(_02113_),
    .A2(_03783_),
    .A3(_03784_),
    .B1(_02332_),
    .B2(\sha256cu.m_out_digest.e_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00245_));
 sky130_fd_sc_hd__nand2_1 _09306_ (.A(_03774_),
    .B(_03775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03785_));
 sky130_fd_sc_hd__or2_1 _09307_ (.A(\sha256cu.m_out_digest.h_in[23] ),
    .B(\sha256cu.m_out_digest.d_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03786_));
 sky130_fd_sc_hd__nand2_1 _09308_ (.A(\sha256cu.m_out_digest.h_in[23] ),
    .B(\sha256cu.m_out_digest.d_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _09309_ (.A(_03786_),
    .B(_03787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03788_));
 sky130_fd_sc_hd__xor2_1 _09310_ (.A(_02851_),
    .B(_03788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03789_));
 sky130_fd_sc_hd__a21boi_1 _09311_ (.A1(_02811_),
    .A2(_03757_),
    .B1_N(_03758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03790_));
 sky130_fd_sc_hd__nor2_1 _09312_ (.A(_03789_),
    .B(_03790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03791_));
 sky130_fd_sc_hd__and2_1 _09313_ (.A(_03789_),
    .B(_03790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03792_));
 sky130_fd_sc_hd__or2_1 _09314_ (.A(_03791_),
    .B(_03792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03793_));
 sky130_fd_sc_hd__inv_2 _09315_ (.A(\sha256cu.K[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03794_));
 sky130_fd_sc_hd__or2_1 _09316_ (.A(\sha256cu.iter_processing.w[23] ),
    .B(_02859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03795_));
 sky130_fd_sc_hd__nand2_1 _09317_ (.A(\sha256cu.iter_processing.w[23] ),
    .B(_02859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _09318_ (.A(_03795_),
    .B(_03796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03797_));
 sky130_fd_sc_hd__xnor2_1 _09319_ (.A(_03794_),
    .B(_03797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03798_));
 sky130_fd_sc_hd__nor2_1 _09320_ (.A(_03793_),
    .B(_03798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03799_));
 sky130_fd_sc_hd__and2_1 _09321_ (.A(_03793_),
    .B(_03798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03800_));
 sky130_fd_sc_hd__nor2_1 _09322_ (.A(_03799_),
    .B(_03800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03801_));
 sky130_fd_sc_hd__o21a_1 _09323_ (.A1(_03762_),
    .A2(_03769_),
    .B1(_03801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03802_));
 sky130_fd_sc_hd__nor3_1 _09324_ (.A(_03762_),
    .B(_03769_),
    .C(_03801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03803_));
 sky130_fd_sc_hd__nor2_1 _09325_ (.A(_03802_),
    .B(_03803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03804_));
 sky130_fd_sc_hd__a21o_1 _09326_ (.A1(\sha256cu.K[22] ),
    .A2(_03767_),
    .B1(_03766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03805_));
 sky130_fd_sc_hd__xnor2_1 _09327_ (.A(_03804_),
    .B(_03805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03806_));
 sky130_fd_sc_hd__and3_1 _09328_ (.A(_03772_),
    .B(_03785_),
    .C(_03806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03807_));
 sky130_fd_sc_hd__a21oi_1 _09329_ (.A1(_03772_),
    .A2(_03785_),
    .B1(_03806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03808_));
 sky130_fd_sc_hd__nor2_1 _09330_ (.A(_03807_),
    .B(_03808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03809_));
 sky130_fd_sc_hd__a21oi_1 _09331_ (.A1(_03777_),
    .A2(_03784_),
    .B1(_03809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03810_));
 sky130_fd_sc_hd__a31o_1 _09332_ (.A1(_03777_),
    .A2(_03784_),
    .A3(_03809_),
    .B1(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03811_));
 sky130_fd_sc_hd__or2_1 _09333_ (.A(\sha256cu.m_out_digest.e_in[23] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03812_));
 sky130_fd_sc_hd__o211a_1 _09334_ (.A1(_03810_),
    .A2(_03811_),
    .B1(_03812_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00246_));
 sky130_fd_sc_hd__or2_1 _09335_ (.A(\sha256cu.m_out_digest.h_in[24] ),
    .B(\sha256cu.m_out_digest.d_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03813_));
 sky130_fd_sc_hd__nand2_1 _09336_ (.A(\sha256cu.m_out_digest.h_in[24] ),
    .B(\sha256cu.m_out_digest.d_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03814_));
 sky130_fd_sc_hd__nand2_1 _09337_ (.A(_03813_),
    .B(_03814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03815_));
 sky130_fd_sc_hd__xor2_1 _09338_ (.A(_02895_),
    .B(_03815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03816_));
 sky130_fd_sc_hd__a21boi_1 _09339_ (.A1(_02851_),
    .A2(_03786_),
    .B1_N(_03787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03817_));
 sky130_fd_sc_hd__or2_1 _09340_ (.A(_03816_),
    .B(_03817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03818_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_03816_),
    .B(_03817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03819_));
 sky130_fd_sc_hd__nand2_1 _09342_ (.A(_03818_),
    .B(_03819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03820_));
 sky130_fd_sc_hd__nor2_1 _09343_ (.A(\sha256cu.iter_processing.w[24] ),
    .B(_02903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03821_));
 sky130_fd_sc_hd__and2_1 _09344_ (.A(\sha256cu.iter_processing.w[24] ),
    .B(_02903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03822_));
 sky130_fd_sc_hd__nor2_1 _09345_ (.A(_03821_),
    .B(_03822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03823_));
 sky130_fd_sc_hd__xnor2_1 _09346_ (.A(\sha256cu.K[24] ),
    .B(_03823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03824_));
 sky130_fd_sc_hd__xor2_1 _09347_ (.A(_03820_),
    .B(_03824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03825_));
 sky130_fd_sc_hd__o21ai_1 _09348_ (.A1(_03791_),
    .A2(_03799_),
    .B1(_03825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03826_));
 sky130_fd_sc_hd__or3_1 _09349_ (.A(_03791_),
    .B(_03799_),
    .C(_03825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03827_));
 sky130_fd_sc_hd__and2_1 _09350_ (.A(_03826_),
    .B(_03827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03828_));
 sky130_fd_sc_hd__o21ai_1 _09351_ (.A1(_03794_),
    .A2(_03797_),
    .B1(_03796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03829_));
 sky130_fd_sc_hd__xor2_1 _09352_ (.A(_03828_),
    .B(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03830_));
 sky130_fd_sc_hd__a21o_1 _09353_ (.A1(_03804_),
    .A2(_03805_),
    .B1(_03802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03831_));
 sky130_fd_sc_hd__nand2_1 _09354_ (.A(_03830_),
    .B(_03831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03832_));
 sky130_fd_sc_hd__or2_1 _09355_ (.A(_03830_),
    .B(_03831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03833_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(_03832_),
    .B(_03833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_1 _09357_ (.A(_03779_),
    .B(_03809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03835_));
 sky130_fd_sc_hd__inv_2 _09358_ (.A(_03782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03836_));
 sky130_fd_sc_hd__inv_2 _09359_ (.A(_03808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03837_));
 sky130_fd_sc_hd__o221a_1 _09360_ (.A1(_03777_),
    .A2(_03807_),
    .B1(_03835_),
    .B2(_03836_),
    .C1(_03837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03838_));
 sky130_fd_sc_hd__o31a_1 _09361_ (.A1(_03725_),
    .A2(_03780_),
    .A3(_03835_),
    .B1(_03838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03839_));
 sky130_fd_sc_hd__or2_1 _09362_ (.A(_03834_),
    .B(_03839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03840_));
 sky130_fd_sc_hd__a21oi_1 _09363_ (.A1(_03834_),
    .A2(_03839_),
    .B1(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03841_));
 sky130_fd_sc_hd__a221o_1 _09364_ (.A1(\sha256cu.m_out_digest.e_in[24] ),
    .A2(_02732_),
    .B1(_03840_),
    .B2(_03841_),
    .C1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00247_));
 sky130_fd_sc_hd__nand2_1 _09365_ (.A(_03828_),
    .B(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03842_));
 sky130_fd_sc_hd__or2_1 _09366_ (.A(\sha256cu.m_out_digest.h_in[25] ),
    .B(\sha256cu.m_out_digest.d_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03843_));
 sky130_fd_sc_hd__nand2_1 _09367_ (.A(\sha256cu.m_out_digest.h_in[25] ),
    .B(\sha256cu.m_out_digest.d_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _09368_ (.A(_03843_),
    .B(_03844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03845_));
 sky130_fd_sc_hd__xor2_1 _09369_ (.A(_02931_),
    .B(_03845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03846_));
 sky130_fd_sc_hd__a21boi_1 _09370_ (.A1(_02895_),
    .A2(_03813_),
    .B1_N(_03814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03847_));
 sky130_fd_sc_hd__nor2_1 _09371_ (.A(_03846_),
    .B(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03848_));
 sky130_fd_sc_hd__and2_1 _09372_ (.A(_03846_),
    .B(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03849_));
 sky130_fd_sc_hd__or2_1 _09373_ (.A(_03848_),
    .B(_03849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03850_));
 sky130_fd_sc_hd__or2_1 _09374_ (.A(\sha256cu.iter_processing.w[25] ),
    .B(_02939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03851_));
 sky130_fd_sc_hd__inv_2 _09375_ (.A(_03851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03852_));
 sky130_fd_sc_hd__and2_1 _09376_ (.A(\sha256cu.iter_processing.w[25] ),
    .B(_02939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03853_));
 sky130_fd_sc_hd__nor2_1 _09377_ (.A(_03852_),
    .B(_03853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03854_));
 sky130_fd_sc_hd__xnor2_1 _09378_ (.A(\sha256cu.K[25] ),
    .B(_03854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03855_));
 sky130_fd_sc_hd__nor2_1 _09379_ (.A(_03850_),
    .B(_03855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03856_));
 sky130_fd_sc_hd__and2_1 _09380_ (.A(_03850_),
    .B(_03855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03857_));
 sky130_fd_sc_hd__nor2_1 _09381_ (.A(_03856_),
    .B(_03857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03858_));
 sky130_fd_sc_hd__o21a_1 _09382_ (.A1(_03820_),
    .A2(_03824_),
    .B1(_03818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03859_));
 sky130_fd_sc_hd__xnor2_1 _09383_ (.A(_03858_),
    .B(_03859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03860_));
 sky130_fd_sc_hd__a21o_1 _09384_ (.A1(\sha256cu.K[24] ),
    .A2(_03823_),
    .B1(_03822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03861_));
 sky130_fd_sc_hd__xnor2_1 _09385_ (.A(_03860_),
    .B(_03861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03862_));
 sky130_fd_sc_hd__and3_1 _09386_ (.A(_03826_),
    .B(_03842_),
    .C(_03862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03863_));
 sky130_fd_sc_hd__a21o_1 _09387_ (.A1(_03826_),
    .A2(_03842_),
    .B1(_03862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03864_));
 sky130_fd_sc_hd__and2b_1 _09388_ (.A_N(_03863_),
    .B(_03864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03865_));
 sky130_fd_sc_hd__and3_1 _09389_ (.A(_03832_),
    .B(_03840_),
    .C(_03865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03866_));
 sky130_fd_sc_hd__a21oi_1 _09390_ (.A1(_03832_),
    .A2(_03840_),
    .B1(_03865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03867_));
 sky130_fd_sc_hd__or2_1 _09391_ (.A(\sha256cu.m_out_digest.e_in[25] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03868_));
 sky130_fd_sc_hd__o311a_1 _09392_ (.A1(_02220_),
    .A2(_03866_),
    .A3(_03867_),
    .B1(_03868_),
    .C1(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00248_));
 sky130_fd_sc_hd__and2_1 _09393_ (.A(_03832_),
    .B(_03864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03869_));
 sky130_fd_sc_hd__or2_1 _09394_ (.A(\sha256cu.m_out_digest.h_in[26] ),
    .B(\sha256cu.m_out_digest.d_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_1 _09395_ (.A(\sha256cu.m_out_digest.h_in[26] ),
    .B(\sha256cu.m_out_digest.d_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03871_));
 sky130_fd_sc_hd__nand2_1 _09396_ (.A(_03870_),
    .B(_03871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03872_));
 sky130_fd_sc_hd__xor2_1 _09397_ (.A(_02964_),
    .B(_03872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03873_));
 sky130_fd_sc_hd__a21boi_1 _09398_ (.A1(_02931_),
    .A2(_03843_),
    .B1_N(_03844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03874_));
 sky130_fd_sc_hd__or2_1 _09399_ (.A(_03873_),
    .B(_03874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03875_));
 sky130_fd_sc_hd__nand2_1 _09400_ (.A(_03873_),
    .B(_03874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _09401_ (.A(_03875_),
    .B(_03876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03877_));
 sky130_fd_sc_hd__nor2_1 _09402_ (.A(\sha256cu.iter_processing.w[26] ),
    .B(_02971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03878_));
 sky130_fd_sc_hd__and2_1 _09403_ (.A(\sha256cu.iter_processing.w[26] ),
    .B(_02971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03879_));
 sky130_fd_sc_hd__nor2_1 _09404_ (.A(_03878_),
    .B(_03879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03880_));
 sky130_fd_sc_hd__xnor2_1 _09405_ (.A(\sha256cu.K[26] ),
    .B(_03880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03881_));
 sky130_fd_sc_hd__xor2_1 _09406_ (.A(_03877_),
    .B(_03881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03882_));
 sky130_fd_sc_hd__o21ai_1 _09407_ (.A1(_03848_),
    .A2(_03856_),
    .B1(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03883_));
 sky130_fd_sc_hd__or3_1 _09408_ (.A(_03848_),
    .B(_03856_),
    .C(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03884_));
 sky130_fd_sc_hd__and2_1 _09409_ (.A(_03883_),
    .B(_03884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03885_));
 sky130_fd_sc_hd__a21o_1 _09410_ (.A1(\sha256cu.K[25] ),
    .A2(_03851_),
    .B1(_03853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03886_));
 sky130_fd_sc_hd__xor2_1 _09411_ (.A(_03885_),
    .B(_03886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03887_));
 sky130_fd_sc_hd__or2b_1 _09412_ (.A(_03859_),
    .B_N(_03858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03888_));
 sky130_fd_sc_hd__a21bo_1 _09413_ (.A1(_03860_),
    .A2(_03861_),
    .B1_N(_03888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03889_));
 sky130_fd_sc_hd__nand2_1 _09414_ (.A(_03887_),
    .B(_03889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03890_));
 sky130_fd_sc_hd__or2_1 _09415_ (.A(_03887_),
    .B(_03889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03891_));
 sky130_fd_sc_hd__and2_1 _09416_ (.A(_03890_),
    .B(_03891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03892_));
 sky130_fd_sc_hd__inv_2 _09417_ (.A(_03892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03893_));
 sky130_fd_sc_hd__a211o_1 _09418_ (.A1(_03840_),
    .A2(_03869_),
    .B1(_03893_),
    .C1(_03863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03894_));
 sky130_fd_sc_hd__or2b_1 _09419_ (.A(_03834_),
    .B_N(_03865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03895_));
 sky130_fd_sc_hd__or2_1 _09420_ (.A(_03863_),
    .B(_03869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03896_));
 sky130_fd_sc_hd__o211ai_1 _09421_ (.A1(_03839_),
    .A2(_03895_),
    .B1(_03896_),
    .C1(_03893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03897_));
 sky130_fd_sc_hd__a32o_1 _09422_ (.A1(_02113_),
    .A2(_03894_),
    .A3(_03897_),
    .B1(_02332_),
    .B2(\sha256cu.m_out_digest.e_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00249_));
 sky130_fd_sc_hd__nand2_1 _09423_ (.A(_03885_),
    .B(_03886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(\sha256cu.m_out_digest.h_in[27] ),
    .B(\sha256cu.m_out_digest.d_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03899_));
 sky130_fd_sc_hd__or2_1 _09425_ (.A(\sha256cu.m_out_digest.h_in[27] ),
    .B(\sha256cu.m_out_digest.d_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03900_));
 sky130_fd_sc_hd__nand2_1 _09426_ (.A(_03899_),
    .B(_03900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03901_));
 sky130_fd_sc_hd__xor2_1 _09427_ (.A(_03001_),
    .B(_03901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03902_));
 sky130_fd_sc_hd__a21boi_1 _09428_ (.A1(_02964_),
    .A2(_03870_),
    .B1_N(_03871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03903_));
 sky130_fd_sc_hd__nor2_1 _09429_ (.A(_03902_),
    .B(_03903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03904_));
 sky130_fd_sc_hd__and2_1 _09430_ (.A(_03902_),
    .B(_03903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03905_));
 sky130_fd_sc_hd__or2_1 _09431_ (.A(_03904_),
    .B(_03905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03906_));
 sky130_fd_sc_hd__or2_1 _09432_ (.A(\sha256cu.iter_processing.w[27] ),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03907_));
 sky130_fd_sc_hd__inv_2 _09433_ (.A(_03907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03908_));
 sky130_fd_sc_hd__and2_1 _09434_ (.A(\sha256cu.iter_processing.w[27] ),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03909_));
 sky130_fd_sc_hd__nor2_1 _09435_ (.A(_03908_),
    .B(_03909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03910_));
 sky130_fd_sc_hd__xnor2_1 _09436_ (.A(\sha256cu.K[27] ),
    .B(_03910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03911_));
 sky130_fd_sc_hd__nor2_1 _09437_ (.A(_03906_),
    .B(_03911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03912_));
 sky130_fd_sc_hd__and2_1 _09438_ (.A(_03906_),
    .B(_03911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03913_));
 sky130_fd_sc_hd__nor2_1 _09439_ (.A(_03912_),
    .B(_03913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03914_));
 sky130_fd_sc_hd__o21a_1 _09440_ (.A1(_03877_),
    .A2(_03881_),
    .B1(_03875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03915_));
 sky130_fd_sc_hd__xnor2_1 _09441_ (.A(_03914_),
    .B(_03915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03916_));
 sky130_fd_sc_hd__a21o_1 _09442_ (.A1(\sha256cu.K[26] ),
    .A2(_03880_),
    .B1(_03879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03917_));
 sky130_fd_sc_hd__xnor2_1 _09443_ (.A(_03916_),
    .B(_03917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03918_));
 sky130_fd_sc_hd__and3_1 _09444_ (.A(_03883_),
    .B(_03898_),
    .C(_03918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03919_));
 sky130_fd_sc_hd__a21oi_1 _09445_ (.A1(_03883_),
    .A2(_03898_),
    .B1(_03918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03920_));
 sky130_fd_sc_hd__nor2_1 _09446_ (.A(_03919_),
    .B(_03920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03921_));
 sky130_fd_sc_hd__and3_1 _09447_ (.A(_03890_),
    .B(_03894_),
    .C(_03921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03922_));
 sky130_fd_sc_hd__a21oi_1 _09448_ (.A1(_03890_),
    .A2(_03894_),
    .B1(_03921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03923_));
 sky130_fd_sc_hd__or2_1 _09449_ (.A(\sha256cu.m_out_digest.e_in[27] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03924_));
 sky130_fd_sc_hd__o311a_1 _09450_ (.A1(_02220_),
    .A2(_03922_),
    .A3(_03923_),
    .B1(_03924_),
    .C1(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00250_));
 sky130_fd_sc_hd__nand2_1 _09451_ (.A(_03892_),
    .B(_03921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03925_));
 sky130_fd_sc_hd__or2_1 _09452_ (.A(_03896_),
    .B(_03925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03926_));
 sky130_fd_sc_hd__o31a_1 _09453_ (.A1(_03839_),
    .A2(_03895_),
    .A3(_03925_),
    .B1(_03926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03927_));
 sky130_fd_sc_hd__o21ba_1 _09454_ (.A1(_03890_),
    .A2(_03919_),
    .B1_N(_03920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03928_));
 sky130_fd_sc_hd__nand2_1 _09455_ (.A(\sha256cu.m_out_digest.h_in[28] ),
    .B(\sha256cu.m_out_digest.d_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03929_));
 sky130_fd_sc_hd__or2_1 _09456_ (.A(\sha256cu.m_out_digest.h_in[28] ),
    .B(\sha256cu.m_out_digest.d_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_1 _09457_ (.A(_03929_),
    .B(_03930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03931_));
 sky130_fd_sc_hd__xor2_1 _09458_ (.A(_03045_),
    .B(_03931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03932_));
 sky130_fd_sc_hd__a21boi_1 _09459_ (.A1(_03001_),
    .A2(_03900_),
    .B1_N(_03899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03933_));
 sky130_fd_sc_hd__nor2_1 _09460_ (.A(_03932_),
    .B(_03933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03934_));
 sky130_fd_sc_hd__and2_1 _09461_ (.A(_03932_),
    .B(_03933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03935_));
 sky130_fd_sc_hd__or2_1 _09462_ (.A(_03934_),
    .B(_03935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03936_));
 sky130_fd_sc_hd__nor2_1 _09463_ (.A(\sha256cu.iter_processing.w[28] ),
    .B(_03052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03937_));
 sky130_fd_sc_hd__and2_1 _09464_ (.A(\sha256cu.iter_processing.w[28] ),
    .B(_03052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03938_));
 sky130_fd_sc_hd__nor2_1 _09465_ (.A(_03937_),
    .B(_03938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03939_));
 sky130_fd_sc_hd__xnor2_1 _09466_ (.A(\sha256cu.K[28] ),
    .B(_03939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03940_));
 sky130_fd_sc_hd__nor2_1 _09467_ (.A(_03936_),
    .B(_03940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03941_));
 sky130_fd_sc_hd__and2_1 _09468_ (.A(_03936_),
    .B(_03940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03942_));
 sky130_fd_sc_hd__nor2_1 _09469_ (.A(_03941_),
    .B(_03942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03943_));
 sky130_fd_sc_hd__o21ai_1 _09470_ (.A1(_03904_),
    .A2(_03912_),
    .B1(_03943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03944_));
 sky130_fd_sc_hd__or3_1 _09471_ (.A(_03904_),
    .B(_03912_),
    .C(_03943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03945_));
 sky130_fd_sc_hd__and2_1 _09472_ (.A(_03944_),
    .B(_03945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03946_));
 sky130_fd_sc_hd__a21o_1 _09473_ (.A1(\sha256cu.K[27] ),
    .A2(_03907_),
    .B1(_03909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03947_));
 sky130_fd_sc_hd__xor2_1 _09474_ (.A(_03946_),
    .B(_03947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03948_));
 sky130_fd_sc_hd__or2b_1 _09475_ (.A(_03915_),
    .B_N(_03914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03949_));
 sky130_fd_sc_hd__a21bo_1 _09476_ (.A1(_03916_),
    .A2(_03917_),
    .B1_N(_03949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03950_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(_03948_),
    .B(_03950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03951_));
 sky130_fd_sc_hd__or2_1 _09478_ (.A(_03948_),
    .B(_03950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03952_));
 sky130_fd_sc_hd__nand2_1 _09479_ (.A(_03951_),
    .B(_03952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03953_));
 sky130_fd_sc_hd__a21o_1 _09480_ (.A1(_03927_),
    .A2(_03928_),
    .B1(_03953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03954_));
 sky130_fd_sc_hd__and3_1 _09481_ (.A(_03927_),
    .B(_03928_),
    .C(_03953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03955_));
 sky130_fd_sc_hd__nor2_1 _09482_ (.A(_02629_),
    .B(_03955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03956_));
 sky130_fd_sc_hd__a221o_1 _09483_ (.A1(\sha256cu.m_out_digest.e_in[28] ),
    .A2(_02732_),
    .B1(_03954_),
    .B2(_03956_),
    .C1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00251_));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(_03946_),
    .B(_03947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03957_));
 sky130_fd_sc_hd__nand2_1 _09485_ (.A(\sha256cu.m_out_digest.h_in[29] ),
    .B(\sha256cu.m_out_digest.d_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03958_));
 sky130_fd_sc_hd__or2_1 _09486_ (.A(\sha256cu.m_out_digest.h_in[29] ),
    .B(\sha256cu.m_out_digest.d_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03959_));
 sky130_fd_sc_hd__nand2_1 _09487_ (.A(_03958_),
    .B(_03959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03960_));
 sky130_fd_sc_hd__xor2_1 _09488_ (.A(_03082_),
    .B(_03960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03961_));
 sky130_fd_sc_hd__a21boi_1 _09489_ (.A1(_03045_),
    .A2(_03930_),
    .B1_N(_03929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03962_));
 sky130_fd_sc_hd__nor2_1 _09490_ (.A(_03961_),
    .B(_03962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03963_));
 sky130_fd_sc_hd__and2_1 _09491_ (.A(_03961_),
    .B(_03962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03964_));
 sky130_fd_sc_hd__or2_1 _09492_ (.A(_03963_),
    .B(_03964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03965_));
 sky130_fd_sc_hd__or2_1 _09493_ (.A(\sha256cu.iter_processing.w[29] ),
    .B(_03089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03966_));
 sky130_fd_sc_hd__nand2_1 _09494_ (.A(\sha256cu.iter_processing.w[29] ),
    .B(_03089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03967_));
 sky130_fd_sc_hd__nand2_1 _09495_ (.A(_03966_),
    .B(_03967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03968_));
 sky130_fd_sc_hd__xnor2_1 _09496_ (.A(_03075_),
    .B(_03968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03969_));
 sky130_fd_sc_hd__nor2_1 _09497_ (.A(_03965_),
    .B(_03969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03970_));
 sky130_fd_sc_hd__and2_1 _09498_ (.A(_03965_),
    .B(_03969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03971_));
 sky130_fd_sc_hd__nor2_1 _09499_ (.A(_03970_),
    .B(_03971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03972_));
 sky130_fd_sc_hd__o21a_1 _09500_ (.A1(_03934_),
    .A2(_03941_),
    .B1(_03972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03973_));
 sky130_fd_sc_hd__nor3_1 _09501_ (.A(_03934_),
    .B(_03941_),
    .C(_03972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03974_));
 sky130_fd_sc_hd__nor2_1 _09502_ (.A(_03973_),
    .B(_03974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03975_));
 sky130_fd_sc_hd__a21o_1 _09503_ (.A1(\sha256cu.K[28] ),
    .A2(_03939_),
    .B1(_03938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03976_));
 sky130_fd_sc_hd__xnor2_1 _09504_ (.A(_03975_),
    .B(_03976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03977_));
 sky130_fd_sc_hd__a21o_1 _09505_ (.A1(_03944_),
    .A2(_03957_),
    .B1(_03977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03978_));
 sky130_fd_sc_hd__inv_2 _09506_ (.A(_03978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03979_));
 sky130_fd_sc_hd__and3_1 _09507_ (.A(_03944_),
    .B(_03957_),
    .C(_03977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03980_));
 sky130_fd_sc_hd__nor2_1 _09508_ (.A(_03979_),
    .B(_03980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03981_));
 sky130_fd_sc_hd__a21oi_1 _09509_ (.A1(_03951_),
    .A2(_03954_),
    .B1(_03981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03982_));
 sky130_fd_sc_hd__a31o_1 _09510_ (.A1(_03951_),
    .A2(_03954_),
    .A3(_03981_),
    .B1(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03983_));
 sky130_fd_sc_hd__o221a_1 _09511_ (.A1(\sha256cu.m_out_digest.e_in[29] ),
    .A2(_02440_),
    .B1(_03982_),
    .B2(_03983_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00252_));
 sky130_fd_sc_hd__and2_1 _09512_ (.A(_03951_),
    .B(_03978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03984_));
 sky130_fd_sc_hd__nor2_1 _09513_ (.A(\sha256cu.m_out_digest.h_in[30] ),
    .B(\sha256cu.m_out_digest.d_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03985_));
 sky130_fd_sc_hd__and2_1 _09514_ (.A(\sha256cu.m_out_digest.h_in[30] ),
    .B(\sha256cu.m_out_digest.d_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03986_));
 sky130_fd_sc_hd__nor2_1 _09515_ (.A(_03985_),
    .B(_03986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03987_));
 sky130_fd_sc_hd__xnor2_1 _09516_ (.A(_03119_),
    .B(_03987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03988_));
 sky130_fd_sc_hd__a21boi_1 _09517_ (.A1(_03082_),
    .A2(_03959_),
    .B1_N(_03958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03989_));
 sky130_fd_sc_hd__or2_1 _09518_ (.A(_03988_),
    .B(_03989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03990_));
 sky130_fd_sc_hd__nand2_1 _09519_ (.A(_03988_),
    .B(_03989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(_03990_),
    .B(_03991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03992_));
 sky130_fd_sc_hd__nor2_1 _09521_ (.A(\sha256cu.iter_processing.w[30] ),
    .B(_03126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03993_));
 sky130_fd_sc_hd__and2_1 _09522_ (.A(\sha256cu.iter_processing.w[30] ),
    .B(_03126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03994_));
 sky130_fd_sc_hd__nor2_1 _09523_ (.A(_03993_),
    .B(_03994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03995_));
 sky130_fd_sc_hd__xnor2_1 _09524_ (.A(\sha256cu.K[30] ),
    .B(_03995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03996_));
 sky130_fd_sc_hd__xor2_1 _09525_ (.A(_03992_),
    .B(_03996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03997_));
 sky130_fd_sc_hd__o21a_1 _09526_ (.A1(_03963_),
    .A2(_03970_),
    .B1(_03997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03998_));
 sky130_fd_sc_hd__nor3_1 _09527_ (.A(_03963_),
    .B(_03970_),
    .C(_03997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03999_));
 sky130_fd_sc_hd__nor2_1 _09528_ (.A(_03998_),
    .B(_03999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04000_));
 sky130_fd_sc_hd__o21ai_1 _09529_ (.A1(_03075_),
    .A2(_03968_),
    .B1(_03967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04001_));
 sky130_fd_sc_hd__xor2_1 _09530_ (.A(_04000_),
    .B(_04001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04002_));
 sky130_fd_sc_hd__a21o_1 _09531_ (.A1(_03975_),
    .A2(_03976_),
    .B1(_03973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04003_));
 sky130_fd_sc_hd__nand2_1 _09532_ (.A(_04002_),
    .B(_04003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04004_));
 sky130_fd_sc_hd__or2_1 _09533_ (.A(_04002_),
    .B(_04003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04005_));
 sky130_fd_sc_hd__nand2_1 _09534_ (.A(_04004_),
    .B(_04005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04006_));
 sky130_fd_sc_hd__a211o_1 _09535_ (.A1(_03954_),
    .A2(_03984_),
    .B1(_04006_),
    .C1(_03980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04007_));
 sky130_fd_sc_hd__a21o_1 _09536_ (.A1(_03954_),
    .A2(_03984_),
    .B1(_03980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04008_));
 sky130_fd_sc_hd__a21oi_1 _09537_ (.A1(_04006_),
    .A2(_04008_),
    .B1(_02069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04009_));
 sky130_fd_sc_hd__and2_1 _09538_ (.A(\sha256cu.m_out_digest.e_in[30] ),
    .B(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04010_));
 sky130_fd_sc_hd__a211o_1 _09539_ (.A1(_04007_),
    .A2(_04009_),
    .B1(_04010_),
    .C1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00253_));
 sky130_fd_sc_hd__a21oi_1 _09540_ (.A1(\sha256cu.K[30] ),
    .A2(_03995_),
    .B1(_03994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04011_));
 sky130_fd_sc_hd__xnor2_1 _09541_ (.A(\sha256cu.m_out_digest.h_in[31] ),
    .B(\sha256cu.m_out_digest.d_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04012_));
 sky130_fd_sc_hd__xnor2_1 _09542_ (.A(_03159_),
    .B(_04012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04013_));
 sky130_fd_sc_hd__xnor2_1 _09543_ (.A(_04011_),
    .B(_04013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04014_));
 sky130_fd_sc_hd__xor2_1 _09544_ (.A(_03157_),
    .B(_04014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04015_));
 sky130_fd_sc_hd__a21oi_1 _09545_ (.A1(_03119_),
    .A2(_03987_),
    .B1(_03986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04016_));
 sky130_fd_sc_hd__xnor2_1 _09546_ (.A(\sha256cu.K[31] ),
    .B(_04016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04017_));
 sky130_fd_sc_hd__a21oi_1 _09547_ (.A1(_04000_),
    .A2(_04001_),
    .B1(_03998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04018_));
 sky130_fd_sc_hd__o21a_1 _09548_ (.A1(_03992_),
    .A2(_03996_),
    .B1(_03990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04019_));
 sky130_fd_sc_hd__xnor2_1 _09549_ (.A(_04018_),
    .B(_04019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04020_));
 sky130_fd_sc_hd__xnor2_1 _09550_ (.A(_04017_),
    .B(_04020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04021_));
 sky130_fd_sc_hd__xnor2_1 _09551_ (.A(_04015_),
    .B(_04021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04022_));
 sky130_fd_sc_hd__and3_1 _09552_ (.A(_04004_),
    .B(_04007_),
    .C(_04022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04023_));
 sky130_fd_sc_hd__a21oi_1 _09553_ (.A1(_04004_),
    .A2(_04007_),
    .B1(_04022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04024_));
 sky130_fd_sc_hd__or2_1 _09554_ (.A(\sha256cu.m_out_digest.e_in[31] ),
    .B(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04025_));
 sky130_fd_sc_hd__o311a_1 _09555_ (.A1(_02220_),
    .A2(_04023_),
    .A3(_04024_),
    .B1(_04025_),
    .C1(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00254_));
 sky130_fd_sc_hd__a22o_1 _09556_ (.A1(\sha256cu.m_out_digest.f_in[0] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00255_));
 sky130_fd_sc_hd__a22o_1 _09557_ (.A1(\sha256cu.m_out_digest.f_in[1] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00256_));
 sky130_fd_sc_hd__o22a_1 _09558_ (.A1(\sha256cu.m_out_digest.f_in[2] ),
    .A2(_03191_),
    .B1(_03190_),
    .B2(\sha256cu.m_out_digest.e_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00257_));
 sky130_fd_sc_hd__buf_4 _09559_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04026_));
 sky130_fd_sc_hd__o22a_1 _09560_ (.A1(\sha256cu.m_out_digest.f_in[3] ),
    .A2(_03191_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00258_));
 sky130_fd_sc_hd__a22o_1 _09561_ (.A1(\sha256cu.m_out_digest.f_in[4] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00259_));
 sky130_fd_sc_hd__a22o_1 _09562_ (.A1(\sha256cu.m_out_digest.f_in[5] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00260_));
 sky130_fd_sc_hd__a22o_1 _09563_ (.A1(\sha256cu.m_out_digest.f_in[6] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00261_));
 sky130_fd_sc_hd__buf_4 _09564_ (.A(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04027_));
 sky130_fd_sc_hd__o22a_1 _09565_ (.A1(\sha256cu.m_out_digest.f_in[7] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00262_));
 sky130_fd_sc_hd__a22o_1 _09566_ (.A1(\sha256cu.m_out_digest.f_in[8] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00263_));
 sky130_fd_sc_hd__a22o_1 _09567_ (.A1(\sha256cu.m_out_digest.f_in[9] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00264_));
 sky130_fd_sc_hd__a22o_1 _09568_ (.A1(\sha256cu.m_out_digest.f_in[10] ),
    .A2(_03559_),
    .B1(_03192_),
    .B2(\sha256cu.m_out_digest.e_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00265_));
 sky130_fd_sc_hd__o22a_1 _09569_ (.A1(\sha256cu.m_out_digest.f_in[11] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00266_));
 sky130_fd_sc_hd__clkbuf_4 _09570_ (.A(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04028_));
 sky130_fd_sc_hd__a22o_1 _09571_ (.A1(\sha256cu.m_out_digest.f_in[12] ),
    .A2(_03559_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00267_));
 sky130_fd_sc_hd__o22a_1 _09572_ (.A1(\sha256cu.m_out_digest.f_in[13] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00268_));
 sky130_fd_sc_hd__o22a_1 _09573_ (.A1(\sha256cu.m_out_digest.f_in[14] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00269_));
 sky130_fd_sc_hd__clkbuf_4 _09574_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04029_));
 sky130_fd_sc_hd__a22o_1 _09575_ (.A1(\sha256cu.m_out_digest.f_in[15] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00270_));
 sky130_fd_sc_hd__o22a_1 _09576_ (.A1(\sha256cu.m_out_digest.f_in[16] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00271_));
 sky130_fd_sc_hd__a22o_1 _09577_ (.A1(\sha256cu.m_out_digest.f_in[17] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00272_));
 sky130_fd_sc_hd__o22a_1 _09578_ (.A1(\sha256cu.m_out_digest.f_in[18] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00273_));
 sky130_fd_sc_hd__a22o_1 _09579_ (.A1(\sha256cu.m_out_digest.f_in[19] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00274_));
 sky130_fd_sc_hd__a22o_1 _09580_ (.A1(\sha256cu.m_out_digest.f_in[20] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00275_));
 sky130_fd_sc_hd__a22o_1 _09581_ (.A1(\sha256cu.m_out_digest.f_in[21] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00276_));
 sky130_fd_sc_hd__a22o_1 _09582_ (.A1(\sha256cu.m_out_digest.f_in[22] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00277_));
 sky130_fd_sc_hd__a22o_1 _09583_ (.A1(\sha256cu.m_out_digest.f_in[23] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00278_));
 sky130_fd_sc_hd__o22a_1 _09584_ (.A1(\sha256cu.m_out_digest.f_in[24] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00279_));
 sky130_fd_sc_hd__o22a_1 _09585_ (.A1(\sha256cu.m_out_digest.f_in[25] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00280_));
 sky130_fd_sc_hd__a22o_1 _09586_ (.A1(\sha256cu.m_out_digest.f_in[26] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00281_));
 sky130_fd_sc_hd__o22a_1 _09587_ (.A1(\sha256cu.m_out_digest.f_in[27] ),
    .A2(_04027_),
    .B1(_04026_),
    .B2(\sha256cu.m_out_digest.e_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00282_));
 sky130_fd_sc_hd__buf_4 _09588_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04030_));
 sky130_fd_sc_hd__o22a_1 _09589_ (.A1(\sha256cu.m_out_digest.f_in[28] ),
    .A2(_04027_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.e_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00283_));
 sky130_fd_sc_hd__a22o_1 _09590_ (.A1(\sha256cu.m_out_digest.f_in[29] ),
    .A2(_04029_),
    .B1(_04028_),
    .B2(\sha256cu.m_out_digest.e_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00284_));
 sky130_fd_sc_hd__buf_4 _09591_ (.A(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04031_));
 sky130_fd_sc_hd__a22o_1 _09592_ (.A1(\sha256cu.m_out_digest.f_in[30] ),
    .A2(_04029_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.e_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00285_));
 sky130_fd_sc_hd__buf_4 _09593_ (.A(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04032_));
 sky130_fd_sc_hd__o22a_1 _09594_ (.A1(\sha256cu.m_out_digest.f_in[31] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.e_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00286_));
 sky130_fd_sc_hd__o22a_1 _09595_ (.A1(\sha256cu.m_out_digest.g_in[0] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00287_));
 sky130_fd_sc_hd__o22a_1 _09596_ (.A1(\sha256cu.m_out_digest.g_in[1] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00288_));
 sky130_fd_sc_hd__buf_4 _09597_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04033_));
 sky130_fd_sc_hd__a22o_1 _09598_ (.A1(\sha256cu.m_out_digest.g_in[2] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00289_));
 sky130_fd_sc_hd__o22a_1 _09599_ (.A1(\sha256cu.m_out_digest.g_in[3] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00290_));
 sky130_fd_sc_hd__a22o_1 _09600_ (.A1(\sha256cu.m_out_digest.g_in[4] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00291_));
 sky130_fd_sc_hd__o22a_1 _09601_ (.A1(\sha256cu.m_out_digest.g_in[5] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00292_));
 sky130_fd_sc_hd__a22o_1 _09602_ (.A1(\sha256cu.m_out_digest.g_in[6] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00293_));
 sky130_fd_sc_hd__o22a_1 _09603_ (.A1(\sha256cu.m_out_digest.g_in[7] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00294_));
 sky130_fd_sc_hd__o22a_1 _09604_ (.A1(\sha256cu.m_out_digest.g_in[8] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00295_));
 sky130_fd_sc_hd__a22o_1 _09605_ (.A1(\sha256cu.m_out_digest.g_in[9] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00296_));
 sky130_fd_sc_hd__a22o_1 _09606_ (.A1(\sha256cu.m_out_digest.g_in[10] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00297_));
 sky130_fd_sc_hd__o22a_1 _09607_ (.A1(\sha256cu.m_out_digest.g_in[11] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00298_));
 sky130_fd_sc_hd__o22a_1 _09608_ (.A1(\sha256cu.m_out_digest.g_in[12] ),
    .A2(_04032_),
    .B1(_04030_),
    .B2(\sha256cu.m_out_digest.f_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00299_));
 sky130_fd_sc_hd__a22o_1 _09609_ (.A1(\sha256cu.m_out_digest.g_in[13] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00300_));
 sky130_fd_sc_hd__clkbuf_4 _09610_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04034_));
 sky130_fd_sc_hd__o22a_1 _09611_ (.A1(\sha256cu.m_out_digest.g_in[14] ),
    .A2(_04032_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00301_));
 sky130_fd_sc_hd__clkbuf_4 _09612_ (.A(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04035_));
 sky130_fd_sc_hd__o22a_1 _09613_ (.A1(\sha256cu.m_out_digest.g_in[15] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00302_));
 sky130_fd_sc_hd__o22a_1 _09614_ (.A1(\sha256cu.m_out_digest.g_in[16] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00303_));
 sky130_fd_sc_hd__o22a_1 _09615_ (.A1(\sha256cu.m_out_digest.g_in[17] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00304_));
 sky130_fd_sc_hd__a22o_1 _09616_ (.A1(\sha256cu.m_out_digest.g_in[18] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00305_));
 sky130_fd_sc_hd__a22o_1 _09617_ (.A1(\sha256cu.m_out_digest.g_in[19] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00306_));
 sky130_fd_sc_hd__a22o_1 _09618_ (.A1(\sha256cu.m_out_digest.g_in[20] ),
    .A2(_04033_),
    .B1(_04031_),
    .B2(\sha256cu.m_out_digest.f_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00307_));
 sky130_fd_sc_hd__buf_4 _09619_ (.A(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04036_));
 sky130_fd_sc_hd__a22o_1 _09620_ (.A1(\sha256cu.m_out_digest.g_in[21] ),
    .A2(_04033_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.f_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00308_));
 sky130_fd_sc_hd__buf_4 _09621_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04037_));
 sky130_fd_sc_hd__a22o_1 _09622_ (.A1(\sha256cu.m_out_digest.g_in[22] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.f_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00309_));
 sky130_fd_sc_hd__o22a_1 _09623_ (.A1(\sha256cu.m_out_digest.g_in[23] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00310_));
 sky130_fd_sc_hd__o22a_1 _09624_ (.A1(\sha256cu.m_out_digest.g_in[24] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00311_));
 sky130_fd_sc_hd__o22a_1 _09625_ (.A1(\sha256cu.m_out_digest.g_in[25] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00312_));
 sky130_fd_sc_hd__o22a_1 _09626_ (.A1(\sha256cu.m_out_digest.g_in[26] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00313_));
 sky130_fd_sc_hd__o22a_1 _09627_ (.A1(\sha256cu.m_out_digest.g_in[27] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00314_));
 sky130_fd_sc_hd__o22a_1 _09628_ (.A1(\sha256cu.m_out_digest.g_in[28] ),
    .A2(_04035_),
    .B1(_04034_),
    .B2(\sha256cu.m_out_digest.f_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00315_));
 sky130_fd_sc_hd__a22o_1 _09629_ (.A1(\sha256cu.m_out_digest.g_in[29] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.f_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00316_));
 sky130_fd_sc_hd__a22o_1 _09630_ (.A1(\sha256cu.m_out_digest.g_in[30] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.f_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00317_));
 sky130_fd_sc_hd__a22o_1 _09631_ (.A1(\sha256cu.m_out_digest.g_in[31] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.f_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00318_));
 sky130_fd_sc_hd__buf_4 _09632_ (.A(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04038_));
 sky130_fd_sc_hd__o22a_1 _09633_ (.A1(\sha256cu.m_out_digest.h_in[0] ),
    .A2(_04035_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00319_));
 sky130_fd_sc_hd__a22o_1 _09634_ (.A1(\sha256cu.m_out_digest.h_in[1] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.g_in[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00320_));
 sky130_fd_sc_hd__a22o_1 _09635_ (.A1(\sha256cu.m_out_digest.h_in[2] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.g_in[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00321_));
 sky130_fd_sc_hd__buf_4 _09636_ (.A(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04039_));
 sky130_fd_sc_hd__o22a_1 _09637_ (.A1(\sha256cu.m_out_digest.h_in[3] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00322_));
 sky130_fd_sc_hd__o22a_1 _09638_ (.A1(\sha256cu.m_out_digest.h_in[4] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00323_));
 sky130_fd_sc_hd__a22o_1 _09639_ (.A1(\sha256cu.m_out_digest.h_in[5] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.g_in[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00324_));
 sky130_fd_sc_hd__a22o_1 _09640_ (.A1(\sha256cu.m_out_digest.h_in[6] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.g_in[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00325_));
 sky130_fd_sc_hd__a22o_1 _09641_ (.A1(\sha256cu.m_out_digest.h_in[7] ),
    .A2(_04037_),
    .B1(_04036_),
    .B2(\sha256cu.m_out_digest.g_in[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00326_));
 sky130_fd_sc_hd__o22a_1 _09642_ (.A1(\sha256cu.m_out_digest.h_in[8] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00327_));
 sky130_fd_sc_hd__clkbuf_4 _09643_ (.A(_02112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04040_));
 sky130_fd_sc_hd__a22o_1 _09644_ (.A1(\sha256cu.m_out_digest.h_in[9] ),
    .A2(_04037_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00328_));
 sky130_fd_sc_hd__o22a_1 _09645_ (.A1(\sha256cu.m_out_digest.h_in[10] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00329_));
 sky130_fd_sc_hd__o22a_1 _09646_ (.A1(\sha256cu.m_out_digest.h_in[11] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00330_));
 sky130_fd_sc_hd__clkbuf_4 _09647_ (.A(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04041_));
 sky130_fd_sc_hd__a22o_1 _09648_ (.A1(\sha256cu.m_out_digest.h_in[12] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00331_));
 sky130_fd_sc_hd__a22o_1 _09649_ (.A1(\sha256cu.m_out_digest.h_in[13] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00332_));
 sky130_fd_sc_hd__o22a_1 _09650_ (.A1(\sha256cu.m_out_digest.h_in[14] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00333_));
 sky130_fd_sc_hd__o22a_1 _09651_ (.A1(\sha256cu.m_out_digest.h_in[15] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00334_));
 sky130_fd_sc_hd__a22o_1 _09652_ (.A1(\sha256cu.m_out_digest.h_in[16] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00335_));
 sky130_fd_sc_hd__a22o_1 _09653_ (.A1(\sha256cu.m_out_digest.h_in[17] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00336_));
 sky130_fd_sc_hd__a22o_1 _09654_ (.A1(\sha256cu.m_out_digest.h_in[18] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00337_));
 sky130_fd_sc_hd__a22o_1 _09655_ (.A1(\sha256cu.m_out_digest.h_in[19] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00338_));
 sky130_fd_sc_hd__a22o_1 _09656_ (.A1(\sha256cu.m_out_digest.h_in[20] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00339_));
 sky130_fd_sc_hd__o22a_1 _09657_ (.A1(\sha256cu.m_out_digest.h_in[21] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00340_));
 sky130_fd_sc_hd__o22a_1 _09658_ (.A1(\sha256cu.m_out_digest.h_in[22] ),
    .A2(_04039_),
    .B1(_04038_),
    .B2(\sha256cu.m_out_digest.g_in[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00341_));
 sky130_fd_sc_hd__o22a_1 _09659_ (.A1(\sha256cu.m_out_digest.h_in[23] ),
    .A2(_04039_),
    .B1(_02478_),
    .B2(\sha256cu.m_out_digest.g_in[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00342_));
 sky130_fd_sc_hd__o22a_1 _09660_ (.A1(\sha256cu.m_out_digest.h_in[24] ),
    .A2(_02369_),
    .B1(_02478_),
    .B2(\sha256cu.m_out_digest.g_in[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00343_));
 sky130_fd_sc_hd__o22a_1 _09661_ (.A1(\sha256cu.m_out_digest.h_in[25] ),
    .A2(_02369_),
    .B1(_02478_),
    .B2(\sha256cu.m_out_digest.g_in[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00344_));
 sky130_fd_sc_hd__a22o_1 _09662_ (.A1(\sha256cu.m_out_digest.h_in[26] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00345_));
 sky130_fd_sc_hd__o22a_1 _09663_ (.A1(\sha256cu.m_out_digest.h_in[27] ),
    .A2(_02369_),
    .B1(_02478_),
    .B2(\sha256cu.m_out_digest.g_in[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00346_));
 sky130_fd_sc_hd__o22a_1 _09664_ (.A1(\sha256cu.m_out_digest.h_in[28] ),
    .A2(_02369_),
    .B1(_02478_),
    .B2(\sha256cu.m_out_digest.g_in[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00347_));
 sky130_fd_sc_hd__a22o_1 _09665_ (.A1(\sha256cu.m_out_digest.h_in[29] ),
    .A2(_04041_),
    .B1(_04040_),
    .B2(\sha256cu.m_out_digest.g_in[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00348_));
 sky130_fd_sc_hd__o22a_1 _09666_ (.A1(\sha256cu.m_out_digest.h_in[30] ),
    .A2(_02369_),
    .B1(_02478_),
    .B2(\sha256cu.m_out_digest.g_in[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00349_));
 sky130_fd_sc_hd__a22o_1 _09667_ (.A1(\sha256cu.m_out_digest.h_in[31] ),
    .A2(_04041_),
    .B1(_02113_),
    .B2(\sha256cu.m_out_digest.g_in[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00350_));
 sky130_fd_sc_hd__or3_1 _09668_ (.A(\sha256cu.msg_scheduler.counter_iteration[5] ),
    .B(\sha256cu.msg_scheduler.counter_iteration[4] ),
    .C(_01565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04042_));
 sky130_fd_sc_hd__buf_6 _09669_ (.A(_04042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_4 _09670_ (.A(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04044_));
 sky130_fd_sc_hd__buf_2 _09671_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_4 _09672_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04046_));
 sky130_fd_sc_hd__or2_1 _09673_ (.A(\sha256cu.iter_processing.w[0] ),
    .B(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04047_));
 sky130_fd_sc_hd__o211a_1 _09674_ (.A1(\sha256cu.msg_scheduler.mreg_14[0] ),
    .A2(_04045_),
    .B1(_04047_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00351_));
 sky130_fd_sc_hd__or2_1 _09675_ (.A(\sha256cu.iter_processing.w[1] ),
    .B(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04048_));
 sky130_fd_sc_hd__o211a_1 _09676_ (.A1(\sha256cu.msg_scheduler.mreg_14[1] ),
    .A2(_04045_),
    .B1(_04048_),
    .C1(_03366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00352_));
 sky130_fd_sc_hd__or2_1 _09677_ (.A(\sha256cu.iter_processing.w[2] ),
    .B(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04049_));
 sky130_fd_sc_hd__buf_2 _09678_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04050_));
 sky130_fd_sc_hd__o211a_1 _09679_ (.A1(\sha256cu.msg_scheduler.mreg_14[2] ),
    .A2(_04045_),
    .B1(_04049_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00353_));
 sky130_fd_sc_hd__or2_1 _09680_ (.A(\sha256cu.iter_processing.w[3] ),
    .B(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04051_));
 sky130_fd_sc_hd__o211a_1 _09681_ (.A1(\sha256cu.msg_scheduler.mreg_14[3] ),
    .A2(_04045_),
    .B1(_04051_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00354_));
 sky130_fd_sc_hd__or2_1 _09682_ (.A(\sha256cu.iter_processing.w[4] ),
    .B(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04052_));
 sky130_fd_sc_hd__o211a_1 _09683_ (.A1(\sha256cu.msg_scheduler.mreg_14[4] ),
    .A2(_04045_),
    .B1(_04052_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00355_));
 sky130_fd_sc_hd__clkbuf_4 _09684_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04053_));
 sky130_fd_sc_hd__clkbuf_2 _09685_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04054_));
 sky130_fd_sc_hd__or2_1 _09686_ (.A(\sha256cu.iter_processing.w[5] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04055_));
 sky130_fd_sc_hd__o211a_1 _09687_ (.A1(\sha256cu.msg_scheduler.mreg_14[5] ),
    .A2(_04045_),
    .B1(_04055_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00356_));
 sky130_fd_sc_hd__or2_1 _09688_ (.A(\sha256cu.iter_processing.w[6] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04056_));
 sky130_fd_sc_hd__o211a_1 _09689_ (.A1(\sha256cu.msg_scheduler.mreg_14[6] ),
    .A2(_04045_),
    .B1(_04056_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00357_));
 sky130_fd_sc_hd__or2_1 _09690_ (.A(\sha256cu.iter_processing.w[7] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04057_));
 sky130_fd_sc_hd__o211a_1 _09691_ (.A1(\sha256cu.msg_scheduler.mreg_14[7] ),
    .A2(_04045_),
    .B1(_04057_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00358_));
 sky130_fd_sc_hd__or2_1 _09692_ (.A(\sha256cu.iter_processing.w[8] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04058_));
 sky130_fd_sc_hd__o211a_1 _09693_ (.A1(\sha256cu.msg_scheduler.mreg_14[8] ),
    .A2(_04045_),
    .B1(_04058_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00359_));
 sky130_fd_sc_hd__or2_1 _09694_ (.A(\sha256cu.iter_processing.w[9] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04059_));
 sky130_fd_sc_hd__o211a_1 _09695_ (.A1(\sha256cu.msg_scheduler.mreg_14[9] ),
    .A2(_04045_),
    .B1(_04059_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00360_));
 sky130_fd_sc_hd__buf_2 _09696_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04060_));
 sky130_fd_sc_hd__or2_1 _09697_ (.A(\sha256cu.iter_processing.w[10] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04061_));
 sky130_fd_sc_hd__o211a_1 _09698_ (.A1(\sha256cu.msg_scheduler.mreg_14[10] ),
    .A2(_04060_),
    .B1(_04061_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00361_));
 sky130_fd_sc_hd__or2_1 _09699_ (.A(\sha256cu.iter_processing.w[11] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04062_));
 sky130_fd_sc_hd__o211a_1 _09700_ (.A1(\sha256cu.msg_scheduler.mreg_14[11] ),
    .A2(_04060_),
    .B1(_04062_),
    .C1(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00362_));
 sky130_fd_sc_hd__or2_1 _09701_ (.A(\sha256cu.iter_processing.w[12] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04063_));
 sky130_fd_sc_hd__buf_2 _09702_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04064_));
 sky130_fd_sc_hd__o211a_1 _09703_ (.A1(\sha256cu.msg_scheduler.mreg_14[12] ),
    .A2(_04060_),
    .B1(_04063_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00363_));
 sky130_fd_sc_hd__or2_1 _09704_ (.A(\sha256cu.iter_processing.w[13] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04065_));
 sky130_fd_sc_hd__o211a_1 _09705_ (.A1(\sha256cu.msg_scheduler.mreg_14[13] ),
    .A2(_04060_),
    .B1(_04065_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00364_));
 sky130_fd_sc_hd__or2_1 _09706_ (.A(\sha256cu.iter_processing.w[14] ),
    .B(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04066_));
 sky130_fd_sc_hd__o211a_1 _09707_ (.A1(\sha256cu.msg_scheduler.mreg_14[14] ),
    .A2(_04060_),
    .B1(_04066_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00365_));
 sky130_fd_sc_hd__clkbuf_2 _09708_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04067_));
 sky130_fd_sc_hd__or2_1 _09709_ (.A(\sha256cu.iter_processing.w[15] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04068_));
 sky130_fd_sc_hd__o211a_1 _09710_ (.A1(\sha256cu.msg_scheduler.mreg_14[15] ),
    .A2(_04060_),
    .B1(_04068_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00366_));
 sky130_fd_sc_hd__or2_1 _09711_ (.A(\sha256cu.iter_processing.w[16] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04069_));
 sky130_fd_sc_hd__o211a_1 _09712_ (.A1(\sha256cu.msg_scheduler.mreg_14[16] ),
    .A2(_04060_),
    .B1(_04069_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00367_));
 sky130_fd_sc_hd__or2_1 _09713_ (.A(\sha256cu.iter_processing.w[17] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04070_));
 sky130_fd_sc_hd__o211a_1 _09714_ (.A1(\sha256cu.msg_scheduler.mreg_14[17] ),
    .A2(_04060_),
    .B1(_04070_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00368_));
 sky130_fd_sc_hd__or2_1 _09715_ (.A(\sha256cu.iter_processing.w[18] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04071_));
 sky130_fd_sc_hd__o211a_1 _09716_ (.A1(\sha256cu.msg_scheduler.mreg_14[18] ),
    .A2(_04060_),
    .B1(_04071_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00369_));
 sky130_fd_sc_hd__or2_1 _09717_ (.A(\sha256cu.iter_processing.w[19] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04072_));
 sky130_fd_sc_hd__o211a_1 _09718_ (.A1(\sha256cu.msg_scheduler.mreg_14[19] ),
    .A2(_04060_),
    .B1(_04072_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00370_));
 sky130_fd_sc_hd__buf_2 _09719_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04073_));
 sky130_fd_sc_hd__or2_1 _09720_ (.A(\sha256cu.iter_processing.w[20] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04074_));
 sky130_fd_sc_hd__o211a_1 _09721_ (.A1(\sha256cu.msg_scheduler.mreg_14[20] ),
    .A2(_04073_),
    .B1(_04074_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00371_));
 sky130_fd_sc_hd__or2_1 _09722_ (.A(\sha256cu.iter_processing.w[21] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04075_));
 sky130_fd_sc_hd__o211a_1 _09723_ (.A1(\sha256cu.msg_scheduler.mreg_14[21] ),
    .A2(_04073_),
    .B1(_04075_),
    .C1(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00372_));
 sky130_fd_sc_hd__or2_1 _09724_ (.A(\sha256cu.iter_processing.w[22] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04076_));
 sky130_fd_sc_hd__buf_2 _09725_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04077_));
 sky130_fd_sc_hd__o211a_1 _09726_ (.A1(\sha256cu.msg_scheduler.mreg_14[22] ),
    .A2(_04073_),
    .B1(_04076_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00373_));
 sky130_fd_sc_hd__or2_1 _09727_ (.A(\sha256cu.iter_processing.w[23] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04078_));
 sky130_fd_sc_hd__o211a_1 _09728_ (.A1(\sha256cu.msg_scheduler.mreg_14[23] ),
    .A2(_04073_),
    .B1(_04078_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00374_));
 sky130_fd_sc_hd__or2_1 _09729_ (.A(\sha256cu.iter_processing.w[24] ),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04079_));
 sky130_fd_sc_hd__o211a_1 _09730_ (.A1(\sha256cu.msg_scheduler.mreg_14[24] ),
    .A2(_04073_),
    .B1(_04079_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00375_));
 sky130_fd_sc_hd__buf_2 _09731_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04080_));
 sky130_fd_sc_hd__or2_1 _09732_ (.A(\sha256cu.iter_processing.w[25] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04081_));
 sky130_fd_sc_hd__o211a_1 _09733_ (.A1(\sha256cu.msg_scheduler.mreg_14[25] ),
    .A2(_04073_),
    .B1(_04081_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00376_));
 sky130_fd_sc_hd__or2_1 _09734_ (.A(\sha256cu.iter_processing.w[26] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04082_));
 sky130_fd_sc_hd__o211a_1 _09735_ (.A1(\sha256cu.msg_scheduler.mreg_14[26] ),
    .A2(_04073_),
    .B1(_04082_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00377_));
 sky130_fd_sc_hd__or2_1 _09736_ (.A(\sha256cu.iter_processing.w[27] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04083_));
 sky130_fd_sc_hd__o211a_1 _09737_ (.A1(\sha256cu.msg_scheduler.mreg_14[27] ),
    .A2(_04073_),
    .B1(_04083_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00378_));
 sky130_fd_sc_hd__or2_1 _09738_ (.A(\sha256cu.iter_processing.w[28] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04084_));
 sky130_fd_sc_hd__o211a_1 _09739_ (.A1(\sha256cu.msg_scheduler.mreg_14[28] ),
    .A2(_04073_),
    .B1(_04084_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00379_));
 sky130_fd_sc_hd__or2_1 _09740_ (.A(\sha256cu.iter_processing.w[29] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04085_));
 sky130_fd_sc_hd__o211a_1 _09741_ (.A1(\sha256cu.msg_scheduler.mreg_14[29] ),
    .A2(_04073_),
    .B1(_04085_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00380_));
 sky130_fd_sc_hd__clkbuf_4 _09742_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04086_));
 sky130_fd_sc_hd__or2_1 _09743_ (.A(\sha256cu.iter_processing.w[30] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04087_));
 sky130_fd_sc_hd__o211a_1 _09744_ (.A1(\sha256cu.msg_scheduler.mreg_14[30] ),
    .A2(_04086_),
    .B1(_04087_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00381_));
 sky130_fd_sc_hd__or2_1 _09745_ (.A(\sha256cu.iter_processing.w[31] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04088_));
 sky130_fd_sc_hd__o211a_1 _09746_ (.A1(\sha256cu.msg_scheduler.mreg_14[31] ),
    .A2(_04086_),
    .B1(_04088_),
    .C1(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00382_));
 sky130_fd_sc_hd__or2_1 _09747_ (.A(\sha256cu.msg_scheduler.mreg_14[0] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04089_));
 sky130_fd_sc_hd__buf_2 _09748_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04090_));
 sky130_fd_sc_hd__o211a_1 _09749_ (.A1(\sha256cu.msg_scheduler.mreg_13[0] ),
    .A2(_04086_),
    .B1(_04089_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00383_));
 sky130_fd_sc_hd__or2_1 _09750_ (.A(\sha256cu.msg_scheduler.mreg_14[1] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04091_));
 sky130_fd_sc_hd__o211a_1 _09751_ (.A1(\sha256cu.msg_scheduler.mreg_13[1] ),
    .A2(_04086_),
    .B1(_04091_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00384_));
 sky130_fd_sc_hd__or2_1 _09752_ (.A(\sha256cu.msg_scheduler.mreg_14[2] ),
    .B(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04092_));
 sky130_fd_sc_hd__o211a_1 _09753_ (.A1(\sha256cu.msg_scheduler.mreg_13[2] ),
    .A2(_04086_),
    .B1(_04092_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00385_));
 sky130_fd_sc_hd__clkbuf_2 _09754_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04093_));
 sky130_fd_sc_hd__or2_1 _09755_ (.A(\sha256cu.msg_scheduler.mreg_14[3] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04094_));
 sky130_fd_sc_hd__o211a_1 _09756_ (.A1(\sha256cu.msg_scheduler.mreg_13[3] ),
    .A2(_04086_),
    .B1(_04094_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00386_));
 sky130_fd_sc_hd__or2_1 _09757_ (.A(\sha256cu.msg_scheduler.mreg_14[4] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04095_));
 sky130_fd_sc_hd__o211a_1 _09758_ (.A1(\sha256cu.msg_scheduler.mreg_13[4] ),
    .A2(_04086_),
    .B1(_04095_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00387_));
 sky130_fd_sc_hd__or2_1 _09759_ (.A(\sha256cu.msg_scheduler.mreg_14[5] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04096_));
 sky130_fd_sc_hd__o211a_1 _09760_ (.A1(\sha256cu.msg_scheduler.mreg_13[5] ),
    .A2(_04086_),
    .B1(_04096_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00388_));
 sky130_fd_sc_hd__or2_1 _09761_ (.A(\sha256cu.msg_scheduler.mreg_14[6] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04097_));
 sky130_fd_sc_hd__o211a_1 _09762_ (.A1(\sha256cu.msg_scheduler.mreg_13[6] ),
    .A2(_04086_),
    .B1(_04097_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00389_));
 sky130_fd_sc_hd__or2_1 _09763_ (.A(\sha256cu.msg_scheduler.mreg_14[7] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04098_));
 sky130_fd_sc_hd__o211a_1 _09764_ (.A1(\sha256cu.msg_scheduler.mreg_13[7] ),
    .A2(_04086_),
    .B1(_04098_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00390_));
 sky130_fd_sc_hd__buf_2 _09765_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04099_));
 sky130_fd_sc_hd__or2_1 _09766_ (.A(\sha256cu.msg_scheduler.mreg_14[8] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04100_));
 sky130_fd_sc_hd__o211a_1 _09767_ (.A1(\sha256cu.msg_scheduler.mreg_13[8] ),
    .A2(_04099_),
    .B1(_04100_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00391_));
 sky130_fd_sc_hd__or2_1 _09768_ (.A(\sha256cu.msg_scheduler.mreg_14[9] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04101_));
 sky130_fd_sc_hd__o211a_1 _09769_ (.A1(\sha256cu.msg_scheduler.mreg_13[9] ),
    .A2(_04099_),
    .B1(_04101_),
    .C1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00392_));
 sky130_fd_sc_hd__or2_1 _09770_ (.A(\sha256cu.msg_scheduler.mreg_14[10] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04102_));
 sky130_fd_sc_hd__buf_2 _09771_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04103_));
 sky130_fd_sc_hd__o211a_1 _09772_ (.A1(\sha256cu.msg_scheduler.mreg_13[10] ),
    .A2(_04099_),
    .B1(_04102_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00393_));
 sky130_fd_sc_hd__or2_1 _09773_ (.A(\sha256cu.msg_scheduler.mreg_14[11] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04104_));
 sky130_fd_sc_hd__o211a_1 _09774_ (.A1(\sha256cu.msg_scheduler.mreg_13[11] ),
    .A2(_04099_),
    .B1(_04104_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00394_));
 sky130_fd_sc_hd__or2_1 _09775_ (.A(\sha256cu.msg_scheduler.mreg_14[12] ),
    .B(_04093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04105_));
 sky130_fd_sc_hd__o211a_1 _09776_ (.A1(\sha256cu.msg_scheduler.mreg_13[12] ),
    .A2(_04099_),
    .B1(_04105_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00395_));
 sky130_fd_sc_hd__clkbuf_2 _09777_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04106_));
 sky130_fd_sc_hd__or2_1 _09778_ (.A(\sha256cu.msg_scheduler.mreg_14[13] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04107_));
 sky130_fd_sc_hd__o211a_1 _09779_ (.A1(\sha256cu.msg_scheduler.mreg_13[13] ),
    .A2(_04099_),
    .B1(_04107_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00396_));
 sky130_fd_sc_hd__or2_1 _09780_ (.A(\sha256cu.msg_scheduler.mreg_14[14] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04108_));
 sky130_fd_sc_hd__o211a_1 _09781_ (.A1(\sha256cu.msg_scheduler.mreg_13[14] ),
    .A2(_04099_),
    .B1(_04108_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00397_));
 sky130_fd_sc_hd__or2_1 _09782_ (.A(\sha256cu.msg_scheduler.mreg_14[15] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04109_));
 sky130_fd_sc_hd__o211a_1 _09783_ (.A1(\sha256cu.msg_scheduler.mreg_13[15] ),
    .A2(_04099_),
    .B1(_04109_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00398_));
 sky130_fd_sc_hd__or2_1 _09784_ (.A(\sha256cu.msg_scheduler.mreg_14[16] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04110_));
 sky130_fd_sc_hd__o211a_1 _09785_ (.A1(\sha256cu.msg_scheduler.mreg_13[16] ),
    .A2(_04099_),
    .B1(_04110_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00399_));
 sky130_fd_sc_hd__or2_1 _09786_ (.A(\sha256cu.msg_scheduler.mreg_14[17] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04111_));
 sky130_fd_sc_hd__o211a_1 _09787_ (.A1(\sha256cu.msg_scheduler.mreg_13[17] ),
    .A2(_04099_),
    .B1(_04111_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00400_));
 sky130_fd_sc_hd__buf_2 _09788_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04112_));
 sky130_fd_sc_hd__or2_1 _09789_ (.A(\sha256cu.msg_scheduler.mreg_14[18] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04113_));
 sky130_fd_sc_hd__o211a_1 _09790_ (.A1(\sha256cu.msg_scheduler.mreg_13[18] ),
    .A2(_04112_),
    .B1(_04113_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00401_));
 sky130_fd_sc_hd__or2_1 _09791_ (.A(\sha256cu.msg_scheduler.mreg_14[19] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04114_));
 sky130_fd_sc_hd__o211a_1 _09792_ (.A1(\sha256cu.msg_scheduler.mreg_13[19] ),
    .A2(_04112_),
    .B1(_04114_),
    .C1(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00402_));
 sky130_fd_sc_hd__or2_1 _09793_ (.A(\sha256cu.msg_scheduler.mreg_14[20] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04115_));
 sky130_fd_sc_hd__buf_4 _09794_ (.A(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04116_));
 sky130_fd_sc_hd__buf_2 _09795_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04117_));
 sky130_fd_sc_hd__o211a_1 _09796_ (.A1(\sha256cu.msg_scheduler.mreg_13[20] ),
    .A2(_04112_),
    .B1(_04115_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00403_));
 sky130_fd_sc_hd__or2_1 _09797_ (.A(\sha256cu.msg_scheduler.mreg_14[21] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04118_));
 sky130_fd_sc_hd__o211a_1 _09798_ (.A1(\sha256cu.msg_scheduler.mreg_13[21] ),
    .A2(_04112_),
    .B1(_04118_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00404_));
 sky130_fd_sc_hd__or2_1 _09799_ (.A(\sha256cu.msg_scheduler.mreg_14[22] ),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04119_));
 sky130_fd_sc_hd__o211a_1 _09800_ (.A1(\sha256cu.msg_scheduler.mreg_13[22] ),
    .A2(_04112_),
    .B1(_04119_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00405_));
 sky130_fd_sc_hd__clkbuf_2 _09801_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04120_));
 sky130_fd_sc_hd__or2_1 _09802_ (.A(\sha256cu.msg_scheduler.mreg_14[23] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04121_));
 sky130_fd_sc_hd__o211a_1 _09803_ (.A1(\sha256cu.msg_scheduler.mreg_13[23] ),
    .A2(_04112_),
    .B1(_04121_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00406_));
 sky130_fd_sc_hd__or2_1 _09804_ (.A(\sha256cu.msg_scheduler.mreg_14[24] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04122_));
 sky130_fd_sc_hd__o211a_1 _09805_ (.A1(\sha256cu.msg_scheduler.mreg_13[24] ),
    .A2(_04112_),
    .B1(_04122_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00407_));
 sky130_fd_sc_hd__or2_1 _09806_ (.A(\sha256cu.msg_scheduler.mreg_14[25] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04123_));
 sky130_fd_sc_hd__o211a_1 _09807_ (.A1(\sha256cu.msg_scheduler.mreg_13[25] ),
    .A2(_04112_),
    .B1(_04123_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00408_));
 sky130_fd_sc_hd__or2_1 _09808_ (.A(\sha256cu.msg_scheduler.mreg_14[26] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04124_));
 sky130_fd_sc_hd__o211a_1 _09809_ (.A1(\sha256cu.msg_scheduler.mreg_13[26] ),
    .A2(_04112_),
    .B1(_04124_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00409_));
 sky130_fd_sc_hd__or2_1 _09810_ (.A(\sha256cu.msg_scheduler.mreg_14[27] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04125_));
 sky130_fd_sc_hd__o211a_1 _09811_ (.A1(\sha256cu.msg_scheduler.mreg_13[27] ),
    .A2(_04112_),
    .B1(_04125_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00410_));
 sky130_fd_sc_hd__buf_2 _09812_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04126_));
 sky130_fd_sc_hd__or2_1 _09813_ (.A(\sha256cu.msg_scheduler.mreg_14[28] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04127_));
 sky130_fd_sc_hd__o211a_1 _09814_ (.A1(\sha256cu.msg_scheduler.mreg_13[28] ),
    .A2(_04126_),
    .B1(_04127_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00411_));
 sky130_fd_sc_hd__or2_1 _09815_ (.A(\sha256cu.msg_scheduler.mreg_14[29] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04128_));
 sky130_fd_sc_hd__o211a_1 _09816_ (.A1(\sha256cu.msg_scheduler.mreg_13[29] ),
    .A2(_04126_),
    .B1(_04128_),
    .C1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00412_));
 sky130_fd_sc_hd__or2_1 _09817_ (.A(\sha256cu.msg_scheduler.mreg_14[30] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04129_));
 sky130_fd_sc_hd__buf_2 _09818_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04130_));
 sky130_fd_sc_hd__o211a_1 _09819_ (.A1(\sha256cu.msg_scheduler.mreg_13[30] ),
    .A2(_04126_),
    .B1(_04129_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00413_));
 sky130_fd_sc_hd__or2_1 _09820_ (.A(\sha256cu.msg_scheduler.mreg_14[31] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04131_));
 sky130_fd_sc_hd__o211a_1 _09821_ (.A1(\sha256cu.msg_scheduler.mreg_13[31] ),
    .A2(_04126_),
    .B1(_04131_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00414_));
 sky130_fd_sc_hd__or2_1 _09822_ (.A(\sha256cu.msg_scheduler.mreg_13[0] ),
    .B(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04132_));
 sky130_fd_sc_hd__o211a_1 _09823_ (.A1(\sha256cu.msg_scheduler.mreg_12[0] ),
    .A2(_04126_),
    .B1(_04132_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00415_));
 sky130_fd_sc_hd__buf_4 _09824_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_2 _09825_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04134_));
 sky130_fd_sc_hd__or2_1 _09826_ (.A(\sha256cu.msg_scheduler.mreg_13[1] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04135_));
 sky130_fd_sc_hd__o211a_1 _09827_ (.A1(\sha256cu.msg_scheduler.mreg_12[1] ),
    .A2(_04126_),
    .B1(_04135_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00416_));
 sky130_fd_sc_hd__or2_1 _09828_ (.A(\sha256cu.msg_scheduler.mreg_13[2] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04136_));
 sky130_fd_sc_hd__o211a_1 _09829_ (.A1(\sha256cu.msg_scheduler.mreg_12[2] ),
    .A2(_04126_),
    .B1(_04136_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00417_));
 sky130_fd_sc_hd__or2_1 _09830_ (.A(\sha256cu.msg_scheduler.mreg_13[3] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04137_));
 sky130_fd_sc_hd__o211a_1 _09831_ (.A1(\sha256cu.msg_scheduler.mreg_12[3] ),
    .A2(_04126_),
    .B1(_04137_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00418_));
 sky130_fd_sc_hd__or2_1 _09832_ (.A(\sha256cu.msg_scheduler.mreg_13[4] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04138_));
 sky130_fd_sc_hd__o211a_1 _09833_ (.A1(\sha256cu.msg_scheduler.mreg_12[4] ),
    .A2(_04126_),
    .B1(_04138_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00419_));
 sky130_fd_sc_hd__or2_1 _09834_ (.A(\sha256cu.msg_scheduler.mreg_13[5] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04139_));
 sky130_fd_sc_hd__o211a_1 _09835_ (.A1(\sha256cu.msg_scheduler.mreg_12[5] ),
    .A2(_04126_),
    .B1(_04139_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00420_));
 sky130_fd_sc_hd__buf_2 _09836_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04140_));
 sky130_fd_sc_hd__or2_1 _09837_ (.A(\sha256cu.msg_scheduler.mreg_13[6] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04141_));
 sky130_fd_sc_hd__o211a_1 _09838_ (.A1(\sha256cu.msg_scheduler.mreg_12[6] ),
    .A2(_04140_),
    .B1(_04141_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00421_));
 sky130_fd_sc_hd__or2_1 _09839_ (.A(\sha256cu.msg_scheduler.mreg_13[7] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04142_));
 sky130_fd_sc_hd__o211a_1 _09840_ (.A1(\sha256cu.msg_scheduler.mreg_12[7] ),
    .A2(_04140_),
    .B1(_04142_),
    .C1(_04130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00422_));
 sky130_fd_sc_hd__or2_1 _09841_ (.A(\sha256cu.msg_scheduler.mreg_13[8] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04143_));
 sky130_fd_sc_hd__buf_2 _09842_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04144_));
 sky130_fd_sc_hd__o211a_1 _09843_ (.A1(\sha256cu.msg_scheduler.mreg_12[8] ),
    .A2(_04140_),
    .B1(_04143_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00423_));
 sky130_fd_sc_hd__or2_1 _09844_ (.A(\sha256cu.msg_scheduler.mreg_13[9] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04145_));
 sky130_fd_sc_hd__o211a_1 _09845_ (.A1(\sha256cu.msg_scheduler.mreg_12[9] ),
    .A2(_04140_),
    .B1(_04145_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00424_));
 sky130_fd_sc_hd__or2_1 _09846_ (.A(\sha256cu.msg_scheduler.mreg_13[10] ),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04146_));
 sky130_fd_sc_hd__o211a_1 _09847_ (.A1(\sha256cu.msg_scheduler.mreg_12[10] ),
    .A2(_04140_),
    .B1(_04146_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00425_));
 sky130_fd_sc_hd__clkbuf_2 _09848_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04147_));
 sky130_fd_sc_hd__or2_1 _09849_ (.A(\sha256cu.msg_scheduler.mreg_13[11] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04148_));
 sky130_fd_sc_hd__o211a_1 _09850_ (.A1(\sha256cu.msg_scheduler.mreg_12[11] ),
    .A2(_04140_),
    .B1(_04148_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00426_));
 sky130_fd_sc_hd__or2_1 _09851_ (.A(\sha256cu.msg_scheduler.mreg_13[12] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04149_));
 sky130_fd_sc_hd__o211a_1 _09852_ (.A1(\sha256cu.msg_scheduler.mreg_12[12] ),
    .A2(_04140_),
    .B1(_04149_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00427_));
 sky130_fd_sc_hd__or2_1 _09853_ (.A(\sha256cu.msg_scheduler.mreg_13[13] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04150_));
 sky130_fd_sc_hd__o211a_1 _09854_ (.A1(\sha256cu.msg_scheduler.mreg_12[13] ),
    .A2(_04140_),
    .B1(_04150_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00428_));
 sky130_fd_sc_hd__or2_1 _09855_ (.A(\sha256cu.msg_scheduler.mreg_13[14] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04151_));
 sky130_fd_sc_hd__o211a_1 _09856_ (.A1(\sha256cu.msg_scheduler.mreg_12[14] ),
    .A2(_04140_),
    .B1(_04151_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00429_));
 sky130_fd_sc_hd__or2_1 _09857_ (.A(\sha256cu.msg_scheduler.mreg_13[15] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04152_));
 sky130_fd_sc_hd__o211a_1 _09858_ (.A1(\sha256cu.msg_scheduler.mreg_12[15] ),
    .A2(_04140_),
    .B1(_04152_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00430_));
 sky130_fd_sc_hd__buf_2 _09859_ (.A(_04044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04153_));
 sky130_fd_sc_hd__or2_1 _09860_ (.A(\sha256cu.msg_scheduler.mreg_13[16] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04154_));
 sky130_fd_sc_hd__o211a_1 _09861_ (.A1(\sha256cu.msg_scheduler.mreg_12[16] ),
    .A2(_04153_),
    .B1(_04154_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00431_));
 sky130_fd_sc_hd__or2_1 _09862_ (.A(\sha256cu.msg_scheduler.mreg_13[17] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04155_));
 sky130_fd_sc_hd__o211a_1 _09863_ (.A1(\sha256cu.msg_scheduler.mreg_12[17] ),
    .A2(_04153_),
    .B1(_04155_),
    .C1(_04144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00432_));
 sky130_fd_sc_hd__or2_1 _09864_ (.A(\sha256cu.msg_scheduler.mreg_13[18] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04156_));
 sky130_fd_sc_hd__buf_2 _09865_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04157_));
 sky130_fd_sc_hd__o211a_1 _09866_ (.A1(\sha256cu.msg_scheduler.mreg_12[18] ),
    .A2(_04153_),
    .B1(_04156_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00433_));
 sky130_fd_sc_hd__or2_1 _09867_ (.A(\sha256cu.msg_scheduler.mreg_13[19] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04158_));
 sky130_fd_sc_hd__o211a_1 _09868_ (.A1(\sha256cu.msg_scheduler.mreg_12[19] ),
    .A2(_04153_),
    .B1(_04158_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00434_));
 sky130_fd_sc_hd__or2_1 _09869_ (.A(\sha256cu.msg_scheduler.mreg_13[20] ),
    .B(_04147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04159_));
 sky130_fd_sc_hd__o211a_1 _09870_ (.A1(\sha256cu.msg_scheduler.mreg_12[20] ),
    .A2(_04153_),
    .B1(_04159_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00435_));
 sky130_fd_sc_hd__clkbuf_2 _09871_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04160_));
 sky130_fd_sc_hd__or2_1 _09872_ (.A(\sha256cu.msg_scheduler.mreg_13[21] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04161_));
 sky130_fd_sc_hd__o211a_1 _09873_ (.A1(\sha256cu.msg_scheduler.mreg_12[21] ),
    .A2(_04153_),
    .B1(_04161_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00436_));
 sky130_fd_sc_hd__or2_1 _09874_ (.A(\sha256cu.msg_scheduler.mreg_13[22] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04162_));
 sky130_fd_sc_hd__o211a_1 _09875_ (.A1(\sha256cu.msg_scheduler.mreg_12[22] ),
    .A2(_04153_),
    .B1(_04162_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00437_));
 sky130_fd_sc_hd__or2_1 _09876_ (.A(\sha256cu.msg_scheduler.mreg_13[23] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04163_));
 sky130_fd_sc_hd__o211a_1 _09877_ (.A1(\sha256cu.msg_scheduler.mreg_12[23] ),
    .A2(_04153_),
    .B1(_04163_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00438_));
 sky130_fd_sc_hd__or2_1 _09878_ (.A(\sha256cu.msg_scheduler.mreg_13[24] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04164_));
 sky130_fd_sc_hd__o211a_1 _09879_ (.A1(\sha256cu.msg_scheduler.mreg_12[24] ),
    .A2(_04153_),
    .B1(_04164_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00439_));
 sky130_fd_sc_hd__or2_1 _09880_ (.A(\sha256cu.msg_scheduler.mreg_13[25] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04165_));
 sky130_fd_sc_hd__o211a_1 _09881_ (.A1(\sha256cu.msg_scheduler.mreg_12[25] ),
    .A2(_04153_),
    .B1(_04165_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00440_));
 sky130_fd_sc_hd__clkbuf_4 _09882_ (.A(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_4 _09883_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04167_));
 sky130_fd_sc_hd__or2_1 _09884_ (.A(\sha256cu.msg_scheduler.mreg_13[26] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04168_));
 sky130_fd_sc_hd__o211a_1 _09885_ (.A1(\sha256cu.msg_scheduler.mreg_12[26] ),
    .A2(_04167_),
    .B1(_04168_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00441_));
 sky130_fd_sc_hd__or2_1 _09886_ (.A(\sha256cu.msg_scheduler.mreg_13[27] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04169_));
 sky130_fd_sc_hd__o211a_1 _09887_ (.A1(\sha256cu.msg_scheduler.mreg_12[27] ),
    .A2(_04167_),
    .B1(_04169_),
    .C1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00442_));
 sky130_fd_sc_hd__or2_1 _09888_ (.A(\sha256cu.msg_scheduler.mreg_13[28] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04170_));
 sky130_fd_sc_hd__buf_6 _09889_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04171_));
 sky130_fd_sc_hd__o211a_1 _09890_ (.A1(\sha256cu.msg_scheduler.mreg_12[28] ),
    .A2(_04167_),
    .B1(_04170_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00443_));
 sky130_fd_sc_hd__or2_1 _09891_ (.A(\sha256cu.msg_scheduler.mreg_13[29] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04172_));
 sky130_fd_sc_hd__o211a_1 _09892_ (.A1(\sha256cu.msg_scheduler.mreg_12[29] ),
    .A2(_04167_),
    .B1(_04172_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00444_));
 sky130_fd_sc_hd__or2_1 _09893_ (.A(\sha256cu.msg_scheduler.mreg_13[30] ),
    .B(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04173_));
 sky130_fd_sc_hd__o211a_1 _09894_ (.A1(\sha256cu.msg_scheduler.mreg_12[30] ),
    .A2(_04167_),
    .B1(_04173_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00445_));
 sky130_fd_sc_hd__buf_2 _09895_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04174_));
 sky130_fd_sc_hd__or2_1 _09896_ (.A(\sha256cu.msg_scheduler.mreg_13[31] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04175_));
 sky130_fd_sc_hd__o211a_1 _09897_ (.A1(\sha256cu.msg_scheduler.mreg_12[31] ),
    .A2(_04167_),
    .B1(_04175_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00446_));
 sky130_fd_sc_hd__and2_1 _09898_ (.A(\sha256cu.msg_scheduler.counter_iteration[0] ),
    .B(\sha256cu.msg_scheduler.temp_case ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04176_));
 sky130_fd_sc_hd__nand2_2 _09899_ (.A(_01564_),
    .B(\sha256cu.iter_processing.padding_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04177_));
 sky130_fd_sc_hd__and3_1 _09900_ (.A(\sha256cu.msg_scheduler.counter_iteration[0] ),
    .B(\sha256cu.msg_scheduler.temp_case ),
    .C(\sha256cu.msg_scheduler.counter_iteration[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04178_));
 sky130_fd_sc_hd__nor2_1 _09901_ (.A(_04177_),
    .B(_04178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04179_));
 sky130_fd_sc_hd__o21a_1 _09902_ (.A1(\sha256cu.msg_scheduler.counter_iteration[1] ),
    .A2(_04176_),
    .B1(_04179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00447_));
 sky130_fd_sc_hd__a21oi_1 _09903_ (.A1(\sha256cu.msg_scheduler.counter_iteration[2] ),
    .A2(_04178_),
    .B1(_04177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04180_));
 sky130_fd_sc_hd__o21a_1 _09904_ (.A1(\sha256cu.msg_scheduler.counter_iteration[2] ),
    .A2(_04178_),
    .B1(_04180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00448_));
 sky130_fd_sc_hd__and3_1 _09905_ (.A(\sha256cu.msg_scheduler.counter_iteration[3] ),
    .B(\sha256cu.msg_scheduler.counter_iteration[2] ),
    .C(_04178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04181_));
 sky130_fd_sc_hd__a21o_1 _09906_ (.A1(\sha256cu.msg_scheduler.counter_iteration[2] ),
    .A2(_04178_),
    .B1(\sha256cu.msg_scheduler.counter_iteration[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04182_));
 sky130_fd_sc_hd__and3b_1 _09907_ (.A_N(_04181_),
    .B(_02007_),
    .C(_04182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _09908_ (.A(_04183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00449_));
 sky130_fd_sc_hd__xnor2_1 _09909_ (.A(\sha256cu.msg_scheduler.counter_iteration[4] ),
    .B(_04181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04184_));
 sky130_fd_sc_hd__nor2_1 _09910_ (.A(_04177_),
    .B(_04184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00450_));
 sky130_fd_sc_hd__and3_1 _09911_ (.A(\sha256cu.msg_scheduler.counter_iteration[5] ),
    .B(\sha256cu.msg_scheduler.counter_iteration[4] ),
    .C(_04181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04185_));
 sky130_fd_sc_hd__a21o_1 _09912_ (.A1(\sha256cu.msg_scheduler.counter_iteration[4] ),
    .A2(_04181_),
    .B1(\sha256cu.msg_scheduler.counter_iteration[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04186_));
 sky130_fd_sc_hd__and3b_1 _09913_ (.A_N(_04185_),
    .B(_04186_),
    .C(_02007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _09914_ (.A(_04187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00451_));
 sky130_fd_sc_hd__buf_2 _09915_ (.A(\sha256cu.counter_iteration[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04188_));
 sky130_fd_sc_hd__or2_1 _09916_ (.A(_04188_),
    .B(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04189_));
 sky130_fd_sc_hd__o211a_1 _09917_ (.A1(\sha256cu.msg_scheduler.counter_iteration[6] ),
    .A2(_01574_),
    .B1(_04189_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00458_));
 sky130_fd_sc_hd__and2b_1 _09918_ (.A_N(_01567_),
    .B(\sha256cu.iter_processing.padding_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04190_));
 sky130_fd_sc_hd__o21a_1 _09919_ (.A1(\sha256cu.msg_scheduler.temp_case ),
    .A2(_04190_),
    .B1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00459_));
 sky130_fd_sc_hd__or2_1 _09920_ (.A(\sha256cu.msg_scheduler.mreg_1[0] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04191_));
 sky130_fd_sc_hd__o211a_1 _09921_ (.A1(\sha256cu.msg_scheduler.mreg_0[0] ),
    .A2(_04167_),
    .B1(_04191_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00460_));
 sky130_fd_sc_hd__or2_1 _09922_ (.A(\sha256cu.msg_scheduler.mreg_1[1] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04192_));
 sky130_fd_sc_hd__o211a_1 _09923_ (.A1(\sha256cu.msg_scheduler.mreg_0[1] ),
    .A2(_04167_),
    .B1(_04192_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00461_));
 sky130_fd_sc_hd__or2_1 _09924_ (.A(\sha256cu.msg_scheduler.mreg_1[2] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04193_));
 sky130_fd_sc_hd__o211a_1 _09925_ (.A1(\sha256cu.msg_scheduler.mreg_0[2] ),
    .A2(_04167_),
    .B1(_04193_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00462_));
 sky130_fd_sc_hd__or2_1 _09926_ (.A(\sha256cu.msg_scheduler.mreg_1[3] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04194_));
 sky130_fd_sc_hd__o211a_1 _09927_ (.A1(\sha256cu.msg_scheduler.mreg_0[3] ),
    .A2(_04167_),
    .B1(_04194_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00463_));
 sky130_fd_sc_hd__clkbuf_4 _09928_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04195_));
 sky130_fd_sc_hd__or2_1 _09929_ (.A(\sha256cu.msg_scheduler.mreg_1[4] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04196_));
 sky130_fd_sc_hd__o211a_1 _09930_ (.A1(\sha256cu.msg_scheduler.mreg_0[4] ),
    .A2(_04195_),
    .B1(_04196_),
    .C1(_04171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00464_));
 sky130_fd_sc_hd__or2_1 _09931_ (.A(\sha256cu.msg_scheduler.mreg_1[5] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_4 _09932_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04198_));
 sky130_fd_sc_hd__o211a_1 _09933_ (.A1(\sha256cu.msg_scheduler.mreg_0[5] ),
    .A2(_04195_),
    .B1(_04197_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00465_));
 sky130_fd_sc_hd__or2_1 _09934_ (.A(\sha256cu.msg_scheduler.mreg_1[6] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04199_));
 sky130_fd_sc_hd__o211a_1 _09935_ (.A1(\sha256cu.msg_scheduler.mreg_0[6] ),
    .A2(_04195_),
    .B1(_04199_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00466_));
 sky130_fd_sc_hd__or2_1 _09936_ (.A(\sha256cu.msg_scheduler.mreg_1[7] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04200_));
 sky130_fd_sc_hd__o211a_1 _09937_ (.A1(\sha256cu.msg_scheduler.mreg_0[7] ),
    .A2(_04195_),
    .B1(_04200_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00467_));
 sky130_fd_sc_hd__or2_1 _09938_ (.A(\sha256cu.msg_scheduler.mreg_1[8] ),
    .B(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04201_));
 sky130_fd_sc_hd__o211a_1 _09939_ (.A1(\sha256cu.msg_scheduler.mreg_0[8] ),
    .A2(_04195_),
    .B1(_04201_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00468_));
 sky130_fd_sc_hd__buf_2 _09940_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04202_));
 sky130_fd_sc_hd__or2_1 _09941_ (.A(\sha256cu.msg_scheduler.mreg_1[9] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04203_));
 sky130_fd_sc_hd__o211a_1 _09942_ (.A1(\sha256cu.msg_scheduler.mreg_0[9] ),
    .A2(_04195_),
    .B1(_04203_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00469_));
 sky130_fd_sc_hd__or2_1 _09943_ (.A(\sha256cu.msg_scheduler.mreg_1[10] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04204_));
 sky130_fd_sc_hd__o211a_1 _09944_ (.A1(\sha256cu.msg_scheduler.mreg_0[10] ),
    .A2(_04195_),
    .B1(_04204_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00470_));
 sky130_fd_sc_hd__or2_1 _09945_ (.A(\sha256cu.msg_scheduler.mreg_1[11] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04205_));
 sky130_fd_sc_hd__o211a_1 _09946_ (.A1(\sha256cu.msg_scheduler.mreg_0[11] ),
    .A2(_04195_),
    .B1(_04205_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00471_));
 sky130_fd_sc_hd__or2_1 _09947_ (.A(\sha256cu.msg_scheduler.mreg_1[12] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04206_));
 sky130_fd_sc_hd__o211a_1 _09948_ (.A1(\sha256cu.msg_scheduler.mreg_0[12] ),
    .A2(_04195_),
    .B1(_04206_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00472_));
 sky130_fd_sc_hd__or2_1 _09949_ (.A(\sha256cu.msg_scheduler.mreg_1[13] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04207_));
 sky130_fd_sc_hd__o211a_1 _09950_ (.A1(\sha256cu.msg_scheduler.mreg_0[13] ),
    .A2(_04195_),
    .B1(_04207_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00473_));
 sky130_fd_sc_hd__clkbuf_4 _09951_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04208_));
 sky130_fd_sc_hd__or2_1 _09952_ (.A(\sha256cu.msg_scheduler.mreg_1[14] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04209_));
 sky130_fd_sc_hd__o211a_1 _09953_ (.A1(\sha256cu.msg_scheduler.mreg_0[14] ),
    .A2(_04208_),
    .B1(_04209_),
    .C1(_04198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00474_));
 sky130_fd_sc_hd__or2_1 _09954_ (.A(\sha256cu.msg_scheduler.mreg_1[15] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_4 _09955_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04211_));
 sky130_fd_sc_hd__o211a_1 _09956_ (.A1(\sha256cu.msg_scheduler.mreg_0[15] ),
    .A2(_04208_),
    .B1(_04210_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00475_));
 sky130_fd_sc_hd__or2_1 _09957_ (.A(\sha256cu.msg_scheduler.mreg_1[16] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04212_));
 sky130_fd_sc_hd__o211a_1 _09958_ (.A1(\sha256cu.msg_scheduler.mreg_0[16] ),
    .A2(_04208_),
    .B1(_04212_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00476_));
 sky130_fd_sc_hd__or2_1 _09959_ (.A(\sha256cu.msg_scheduler.mreg_1[17] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04213_));
 sky130_fd_sc_hd__o211a_1 _09960_ (.A1(\sha256cu.msg_scheduler.mreg_0[17] ),
    .A2(_04208_),
    .B1(_04213_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00477_));
 sky130_fd_sc_hd__or2_1 _09961_ (.A(\sha256cu.msg_scheduler.mreg_1[18] ),
    .B(_04202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04214_));
 sky130_fd_sc_hd__o211a_1 _09962_ (.A1(\sha256cu.msg_scheduler.mreg_0[18] ),
    .A2(_04208_),
    .B1(_04214_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00478_));
 sky130_fd_sc_hd__clkbuf_2 _09963_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04215_));
 sky130_fd_sc_hd__or2_1 _09964_ (.A(\sha256cu.msg_scheduler.mreg_1[19] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04216_));
 sky130_fd_sc_hd__o211a_1 _09965_ (.A1(\sha256cu.msg_scheduler.mreg_0[19] ),
    .A2(_04208_),
    .B1(_04216_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00479_));
 sky130_fd_sc_hd__or2_1 _09966_ (.A(\sha256cu.msg_scheduler.mreg_1[20] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04217_));
 sky130_fd_sc_hd__o211a_1 _09967_ (.A1(\sha256cu.msg_scheduler.mreg_0[20] ),
    .A2(_04208_),
    .B1(_04217_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00480_));
 sky130_fd_sc_hd__or2_1 _09968_ (.A(\sha256cu.msg_scheduler.mreg_1[21] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04218_));
 sky130_fd_sc_hd__o211a_1 _09969_ (.A1(\sha256cu.msg_scheduler.mreg_0[21] ),
    .A2(_04208_),
    .B1(_04218_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00481_));
 sky130_fd_sc_hd__or2_1 _09970_ (.A(\sha256cu.msg_scheduler.mreg_1[22] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04219_));
 sky130_fd_sc_hd__o211a_1 _09971_ (.A1(\sha256cu.msg_scheduler.mreg_0[22] ),
    .A2(_04208_),
    .B1(_04219_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00482_));
 sky130_fd_sc_hd__or2_1 _09972_ (.A(\sha256cu.msg_scheduler.mreg_1[23] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04220_));
 sky130_fd_sc_hd__o211a_1 _09973_ (.A1(\sha256cu.msg_scheduler.mreg_0[23] ),
    .A2(_04208_),
    .B1(_04220_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00483_));
 sky130_fd_sc_hd__clkbuf_4 _09974_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04221_));
 sky130_fd_sc_hd__or2_1 _09975_ (.A(\sha256cu.msg_scheduler.mreg_1[24] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04222_));
 sky130_fd_sc_hd__o211a_1 _09976_ (.A1(\sha256cu.msg_scheduler.mreg_0[24] ),
    .A2(_04221_),
    .B1(_04222_),
    .C1(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00484_));
 sky130_fd_sc_hd__or2_1 _09977_ (.A(\sha256cu.msg_scheduler.mreg_1[25] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04223_));
 sky130_fd_sc_hd__buf_2 _09978_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04224_));
 sky130_fd_sc_hd__o211a_1 _09979_ (.A1(\sha256cu.msg_scheduler.mreg_0[25] ),
    .A2(_04221_),
    .B1(_04223_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00485_));
 sky130_fd_sc_hd__or2_1 _09980_ (.A(\sha256cu.msg_scheduler.mreg_1[26] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04225_));
 sky130_fd_sc_hd__o211a_1 _09981_ (.A1(\sha256cu.msg_scheduler.mreg_0[26] ),
    .A2(_04221_),
    .B1(_04225_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00486_));
 sky130_fd_sc_hd__or2_1 _09982_ (.A(\sha256cu.msg_scheduler.mreg_1[27] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04226_));
 sky130_fd_sc_hd__o211a_1 _09983_ (.A1(\sha256cu.msg_scheduler.mreg_0[27] ),
    .A2(_04221_),
    .B1(_04226_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00487_));
 sky130_fd_sc_hd__or2_1 _09984_ (.A(\sha256cu.msg_scheduler.mreg_1[28] ),
    .B(_04215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04227_));
 sky130_fd_sc_hd__o211a_1 _09985_ (.A1(\sha256cu.msg_scheduler.mreg_0[28] ),
    .A2(_04221_),
    .B1(_04227_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00488_));
 sky130_fd_sc_hd__clkbuf_2 _09986_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04228_));
 sky130_fd_sc_hd__or2_1 _09987_ (.A(\sha256cu.msg_scheduler.mreg_1[29] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04229_));
 sky130_fd_sc_hd__o211a_1 _09988_ (.A1(\sha256cu.msg_scheduler.mreg_0[29] ),
    .A2(_04221_),
    .B1(_04229_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00489_));
 sky130_fd_sc_hd__or2_1 _09989_ (.A(\sha256cu.msg_scheduler.mreg_1[30] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04230_));
 sky130_fd_sc_hd__o211a_1 _09990_ (.A1(\sha256cu.msg_scheduler.mreg_0[30] ),
    .A2(_04221_),
    .B1(_04230_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00490_));
 sky130_fd_sc_hd__or2_1 _09991_ (.A(\sha256cu.msg_scheduler.mreg_1[31] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04231_));
 sky130_fd_sc_hd__o211a_1 _09992_ (.A1(\sha256cu.msg_scheduler.mreg_0[31] ),
    .A2(_04221_),
    .B1(_04231_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00491_));
 sky130_fd_sc_hd__or2_1 _09993_ (.A(\sha256cu.msg_scheduler.mreg_2[0] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04232_));
 sky130_fd_sc_hd__o211a_1 _09994_ (.A1(\sha256cu.msg_scheduler.mreg_1[0] ),
    .A2(_04221_),
    .B1(_04232_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00492_));
 sky130_fd_sc_hd__or2_1 _09995_ (.A(\sha256cu.msg_scheduler.mreg_2[1] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04233_));
 sky130_fd_sc_hd__o211a_1 _09996_ (.A1(\sha256cu.msg_scheduler.mreg_1[1] ),
    .A2(_04221_),
    .B1(_04233_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00493_));
 sky130_fd_sc_hd__buf_2 _09997_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04234_));
 sky130_fd_sc_hd__or2_1 _09998_ (.A(\sha256cu.msg_scheduler.mreg_2[2] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04235_));
 sky130_fd_sc_hd__o211a_1 _09999_ (.A1(\sha256cu.msg_scheduler.mreg_1[2] ),
    .A2(_04234_),
    .B1(_04235_),
    .C1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00494_));
 sky130_fd_sc_hd__or2_1 _10000_ (.A(\sha256cu.msg_scheduler.mreg_2[3] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04236_));
 sky130_fd_sc_hd__buf_2 _10001_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04237_));
 sky130_fd_sc_hd__o211a_1 _10002_ (.A1(\sha256cu.msg_scheduler.mreg_1[3] ),
    .A2(_04234_),
    .B1(_04236_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00495_));
 sky130_fd_sc_hd__or2_1 _10003_ (.A(\sha256cu.msg_scheduler.mreg_2[4] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04238_));
 sky130_fd_sc_hd__o211a_1 _10004_ (.A1(\sha256cu.msg_scheduler.mreg_1[4] ),
    .A2(_04234_),
    .B1(_04238_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00496_));
 sky130_fd_sc_hd__or2_1 _10005_ (.A(\sha256cu.msg_scheduler.mreg_2[5] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04239_));
 sky130_fd_sc_hd__o211a_1 _10006_ (.A1(\sha256cu.msg_scheduler.mreg_1[5] ),
    .A2(_04234_),
    .B1(_04239_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00497_));
 sky130_fd_sc_hd__or2_1 _10007_ (.A(\sha256cu.msg_scheduler.mreg_2[6] ),
    .B(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04240_));
 sky130_fd_sc_hd__o211a_1 _10008_ (.A1(\sha256cu.msg_scheduler.mreg_1[6] ),
    .A2(_04234_),
    .B1(_04240_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00498_));
 sky130_fd_sc_hd__clkbuf_2 _10009_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04241_));
 sky130_fd_sc_hd__or2_1 _10010_ (.A(\sha256cu.msg_scheduler.mreg_2[7] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04242_));
 sky130_fd_sc_hd__o211a_1 _10011_ (.A1(\sha256cu.msg_scheduler.mreg_1[7] ),
    .A2(_04234_),
    .B1(_04242_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00499_));
 sky130_fd_sc_hd__or2_1 _10012_ (.A(\sha256cu.msg_scheduler.mreg_2[8] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04243_));
 sky130_fd_sc_hd__o211a_1 _10013_ (.A1(\sha256cu.msg_scheduler.mreg_1[8] ),
    .A2(_04234_),
    .B1(_04243_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00500_));
 sky130_fd_sc_hd__or2_1 _10014_ (.A(\sha256cu.msg_scheduler.mreg_2[9] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04244_));
 sky130_fd_sc_hd__o211a_1 _10015_ (.A1(\sha256cu.msg_scheduler.mreg_1[9] ),
    .A2(_04234_),
    .B1(_04244_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00501_));
 sky130_fd_sc_hd__or2_1 _10016_ (.A(\sha256cu.msg_scheduler.mreg_2[10] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04245_));
 sky130_fd_sc_hd__o211a_1 _10017_ (.A1(\sha256cu.msg_scheduler.mreg_1[10] ),
    .A2(_04234_),
    .B1(_04245_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00502_));
 sky130_fd_sc_hd__or2_1 _10018_ (.A(\sha256cu.msg_scheduler.mreg_2[11] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04246_));
 sky130_fd_sc_hd__o211a_1 _10019_ (.A1(\sha256cu.msg_scheduler.mreg_1[11] ),
    .A2(_04234_),
    .B1(_04246_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00503_));
 sky130_fd_sc_hd__buf_2 _10020_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04247_));
 sky130_fd_sc_hd__or2_1 _10021_ (.A(\sha256cu.msg_scheduler.mreg_2[12] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04248_));
 sky130_fd_sc_hd__o211a_1 _10022_ (.A1(\sha256cu.msg_scheduler.mreg_1[12] ),
    .A2(_04247_),
    .B1(_04248_),
    .C1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00504_));
 sky130_fd_sc_hd__or2_1 _10023_ (.A(\sha256cu.msg_scheduler.mreg_2[13] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04249_));
 sky130_fd_sc_hd__buf_2 _10024_ (.A(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04250_));
 sky130_fd_sc_hd__o211a_1 _10025_ (.A1(\sha256cu.msg_scheduler.mreg_1[13] ),
    .A2(_04247_),
    .B1(_04249_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00505_));
 sky130_fd_sc_hd__or2_1 _10026_ (.A(\sha256cu.msg_scheduler.mreg_2[14] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04251_));
 sky130_fd_sc_hd__o211a_1 _10027_ (.A1(\sha256cu.msg_scheduler.mreg_1[14] ),
    .A2(_04247_),
    .B1(_04251_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00506_));
 sky130_fd_sc_hd__or2_1 _10028_ (.A(\sha256cu.msg_scheduler.mreg_2[15] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04252_));
 sky130_fd_sc_hd__o211a_1 _10029_ (.A1(\sha256cu.msg_scheduler.mreg_1[15] ),
    .A2(_04247_),
    .B1(_04252_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00507_));
 sky130_fd_sc_hd__or2_1 _10030_ (.A(\sha256cu.msg_scheduler.mreg_2[16] ),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04253_));
 sky130_fd_sc_hd__o211a_1 _10031_ (.A1(\sha256cu.msg_scheduler.mreg_1[16] ),
    .A2(_04247_),
    .B1(_04253_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00508_));
 sky130_fd_sc_hd__clkbuf_2 _10032_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04254_));
 sky130_fd_sc_hd__or2_1 _10033_ (.A(\sha256cu.msg_scheduler.mreg_2[17] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04255_));
 sky130_fd_sc_hd__o211a_1 _10034_ (.A1(\sha256cu.msg_scheduler.mreg_1[17] ),
    .A2(_04247_),
    .B1(_04255_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00509_));
 sky130_fd_sc_hd__or2_1 _10035_ (.A(\sha256cu.msg_scheduler.mreg_2[18] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04256_));
 sky130_fd_sc_hd__o211a_1 _10036_ (.A1(\sha256cu.msg_scheduler.mreg_1[18] ),
    .A2(_04247_),
    .B1(_04256_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00510_));
 sky130_fd_sc_hd__or2_1 _10037_ (.A(\sha256cu.msg_scheduler.mreg_2[19] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04257_));
 sky130_fd_sc_hd__o211a_1 _10038_ (.A1(\sha256cu.msg_scheduler.mreg_1[19] ),
    .A2(_04247_),
    .B1(_04257_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00511_));
 sky130_fd_sc_hd__or2_1 _10039_ (.A(\sha256cu.msg_scheduler.mreg_2[20] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04258_));
 sky130_fd_sc_hd__o211a_1 _10040_ (.A1(\sha256cu.msg_scheduler.mreg_1[20] ),
    .A2(_04247_),
    .B1(_04258_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00512_));
 sky130_fd_sc_hd__or2_1 _10041_ (.A(\sha256cu.msg_scheduler.mreg_2[21] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04259_));
 sky130_fd_sc_hd__o211a_1 _10042_ (.A1(\sha256cu.msg_scheduler.mreg_1[21] ),
    .A2(_04247_),
    .B1(_04259_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00513_));
 sky130_fd_sc_hd__buf_2 _10043_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04260_));
 sky130_fd_sc_hd__or2_1 _10044_ (.A(\sha256cu.msg_scheduler.mreg_2[22] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04261_));
 sky130_fd_sc_hd__o211a_1 _10045_ (.A1(\sha256cu.msg_scheduler.mreg_1[22] ),
    .A2(_04260_),
    .B1(_04261_),
    .C1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00514_));
 sky130_fd_sc_hd__or2_1 _10046_ (.A(\sha256cu.msg_scheduler.mreg_2[23] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04262_));
 sky130_fd_sc_hd__buf_2 _10047_ (.A(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04263_));
 sky130_fd_sc_hd__buf_2 _10048_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04264_));
 sky130_fd_sc_hd__o211a_1 _10049_ (.A1(\sha256cu.msg_scheduler.mreg_1[23] ),
    .A2(_04260_),
    .B1(_04262_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00515_));
 sky130_fd_sc_hd__or2_1 _10050_ (.A(\sha256cu.msg_scheduler.mreg_2[24] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04265_));
 sky130_fd_sc_hd__o211a_1 _10051_ (.A1(\sha256cu.msg_scheduler.mreg_1[24] ),
    .A2(_04260_),
    .B1(_04265_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00516_));
 sky130_fd_sc_hd__or2_1 _10052_ (.A(\sha256cu.msg_scheduler.mreg_2[25] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04266_));
 sky130_fd_sc_hd__o211a_1 _10053_ (.A1(\sha256cu.msg_scheduler.mreg_1[25] ),
    .A2(_04260_),
    .B1(_04266_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00517_));
 sky130_fd_sc_hd__or2_1 _10054_ (.A(\sha256cu.msg_scheduler.mreg_2[26] ),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04267_));
 sky130_fd_sc_hd__o211a_1 _10055_ (.A1(\sha256cu.msg_scheduler.mreg_1[26] ),
    .A2(_04260_),
    .B1(_04267_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00518_));
 sky130_fd_sc_hd__clkbuf_2 _10056_ (.A(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04268_));
 sky130_fd_sc_hd__or2_1 _10057_ (.A(\sha256cu.msg_scheduler.mreg_2[27] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04269_));
 sky130_fd_sc_hd__o211a_1 _10058_ (.A1(\sha256cu.msg_scheduler.mreg_1[27] ),
    .A2(_04260_),
    .B1(_04269_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00519_));
 sky130_fd_sc_hd__or2_1 _10059_ (.A(\sha256cu.msg_scheduler.mreg_2[28] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04270_));
 sky130_fd_sc_hd__o211a_1 _10060_ (.A1(\sha256cu.msg_scheduler.mreg_1[28] ),
    .A2(_04260_),
    .B1(_04270_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00520_));
 sky130_fd_sc_hd__or2_1 _10061_ (.A(\sha256cu.msg_scheduler.mreg_2[29] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04271_));
 sky130_fd_sc_hd__o211a_1 _10062_ (.A1(\sha256cu.msg_scheduler.mreg_1[29] ),
    .A2(_04260_),
    .B1(_04271_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00521_));
 sky130_fd_sc_hd__or2_1 _10063_ (.A(\sha256cu.msg_scheduler.mreg_2[30] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04272_));
 sky130_fd_sc_hd__o211a_1 _10064_ (.A1(\sha256cu.msg_scheduler.mreg_1[30] ),
    .A2(_04260_),
    .B1(_04272_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00522_));
 sky130_fd_sc_hd__or2_1 _10065_ (.A(\sha256cu.msg_scheduler.mreg_2[31] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04273_));
 sky130_fd_sc_hd__o211a_1 _10066_ (.A1(\sha256cu.msg_scheduler.mreg_1[31] ),
    .A2(_04260_),
    .B1(_04273_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00523_));
 sky130_fd_sc_hd__clkbuf_4 _10067_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04274_));
 sky130_fd_sc_hd__or2_1 _10068_ (.A(\sha256cu.msg_scheduler.mreg_3[0] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04275_));
 sky130_fd_sc_hd__o211a_1 _10069_ (.A1(\sha256cu.msg_scheduler.mreg_2[0] ),
    .A2(_04274_),
    .B1(_04275_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00524_));
 sky130_fd_sc_hd__or2_1 _10070_ (.A(\sha256cu.msg_scheduler.mreg_3[1] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04276_));
 sky130_fd_sc_hd__buf_2 _10071_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04277_));
 sky130_fd_sc_hd__o211a_1 _10072_ (.A1(\sha256cu.msg_scheduler.mreg_2[1] ),
    .A2(_04274_),
    .B1(_04276_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00525_));
 sky130_fd_sc_hd__or2_1 _10073_ (.A(\sha256cu.msg_scheduler.mreg_3[2] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04278_));
 sky130_fd_sc_hd__o211a_1 _10074_ (.A1(\sha256cu.msg_scheduler.mreg_2[2] ),
    .A2(_04274_),
    .B1(_04278_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00526_));
 sky130_fd_sc_hd__or2_1 _10075_ (.A(\sha256cu.msg_scheduler.mreg_3[3] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04279_));
 sky130_fd_sc_hd__o211a_1 _10076_ (.A1(\sha256cu.msg_scheduler.mreg_2[3] ),
    .A2(_04274_),
    .B1(_04279_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00527_));
 sky130_fd_sc_hd__or2_1 _10077_ (.A(\sha256cu.msg_scheduler.mreg_3[4] ),
    .B(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04280_));
 sky130_fd_sc_hd__o211a_1 _10078_ (.A1(\sha256cu.msg_scheduler.mreg_2[4] ),
    .A2(_04274_),
    .B1(_04280_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00528_));
 sky130_fd_sc_hd__clkbuf_4 _10079_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_2 _10080_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04282_));
 sky130_fd_sc_hd__or2_1 _10081_ (.A(\sha256cu.msg_scheduler.mreg_3[5] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04283_));
 sky130_fd_sc_hd__o211a_1 _10082_ (.A1(\sha256cu.msg_scheduler.mreg_2[5] ),
    .A2(_04274_),
    .B1(_04283_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00529_));
 sky130_fd_sc_hd__or2_1 _10083_ (.A(\sha256cu.msg_scheduler.mreg_3[6] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04284_));
 sky130_fd_sc_hd__o211a_1 _10084_ (.A1(\sha256cu.msg_scheduler.mreg_2[6] ),
    .A2(_04274_),
    .B1(_04284_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00530_));
 sky130_fd_sc_hd__or2_1 _10085_ (.A(\sha256cu.msg_scheduler.mreg_3[7] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04285_));
 sky130_fd_sc_hd__o211a_1 _10086_ (.A1(\sha256cu.msg_scheduler.mreg_2[7] ),
    .A2(_04274_),
    .B1(_04285_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00531_));
 sky130_fd_sc_hd__or2_1 _10087_ (.A(\sha256cu.msg_scheduler.mreg_3[8] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04286_));
 sky130_fd_sc_hd__o211a_1 _10088_ (.A1(\sha256cu.msg_scheduler.mreg_2[8] ),
    .A2(_04274_),
    .B1(_04286_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00532_));
 sky130_fd_sc_hd__or2_1 _10089_ (.A(\sha256cu.msg_scheduler.mreg_3[9] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04287_));
 sky130_fd_sc_hd__o211a_1 _10090_ (.A1(\sha256cu.msg_scheduler.mreg_2[9] ),
    .A2(_04274_),
    .B1(_04287_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00533_));
 sky130_fd_sc_hd__buf_2 _10091_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04288_));
 sky130_fd_sc_hd__or2_1 _10092_ (.A(\sha256cu.msg_scheduler.mreg_3[10] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04289_));
 sky130_fd_sc_hd__o211a_1 _10093_ (.A1(\sha256cu.msg_scheduler.mreg_2[10] ),
    .A2(_04288_),
    .B1(_04289_),
    .C1(_04277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00534_));
 sky130_fd_sc_hd__or2_1 _10094_ (.A(\sha256cu.msg_scheduler.mreg_3[11] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04290_));
 sky130_fd_sc_hd__buf_2 _10095_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04291_));
 sky130_fd_sc_hd__o211a_1 _10096_ (.A1(\sha256cu.msg_scheduler.mreg_2[11] ),
    .A2(_04288_),
    .B1(_04290_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00535_));
 sky130_fd_sc_hd__or2_1 _10097_ (.A(\sha256cu.msg_scheduler.mreg_3[12] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04292_));
 sky130_fd_sc_hd__o211a_1 _10098_ (.A1(\sha256cu.msg_scheduler.mreg_2[12] ),
    .A2(_04288_),
    .B1(_04292_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00536_));
 sky130_fd_sc_hd__or2_1 _10099_ (.A(\sha256cu.msg_scheduler.mreg_3[13] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04293_));
 sky130_fd_sc_hd__o211a_1 _10100_ (.A1(\sha256cu.msg_scheduler.mreg_2[13] ),
    .A2(_04288_),
    .B1(_04293_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00537_));
 sky130_fd_sc_hd__or2_1 _10101_ (.A(\sha256cu.msg_scheduler.mreg_3[14] ),
    .B(_04282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04294_));
 sky130_fd_sc_hd__o211a_1 _10102_ (.A1(\sha256cu.msg_scheduler.mreg_2[14] ),
    .A2(_04288_),
    .B1(_04294_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00538_));
 sky130_fd_sc_hd__clkbuf_2 _10103_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04295_));
 sky130_fd_sc_hd__or2_1 _10104_ (.A(\sha256cu.msg_scheduler.mreg_3[15] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04296_));
 sky130_fd_sc_hd__o211a_1 _10105_ (.A1(\sha256cu.msg_scheduler.mreg_2[15] ),
    .A2(_04288_),
    .B1(_04296_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00539_));
 sky130_fd_sc_hd__or2_1 _10106_ (.A(\sha256cu.msg_scheduler.mreg_3[16] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04297_));
 sky130_fd_sc_hd__o211a_1 _10107_ (.A1(\sha256cu.msg_scheduler.mreg_2[16] ),
    .A2(_04288_),
    .B1(_04297_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00540_));
 sky130_fd_sc_hd__or2_1 _10108_ (.A(\sha256cu.msg_scheduler.mreg_3[17] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04298_));
 sky130_fd_sc_hd__o211a_1 _10109_ (.A1(\sha256cu.msg_scheduler.mreg_2[17] ),
    .A2(_04288_),
    .B1(_04298_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00541_));
 sky130_fd_sc_hd__or2_1 _10110_ (.A(\sha256cu.msg_scheduler.mreg_3[18] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04299_));
 sky130_fd_sc_hd__o211a_1 _10111_ (.A1(\sha256cu.msg_scheduler.mreg_2[18] ),
    .A2(_04288_),
    .B1(_04299_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00542_));
 sky130_fd_sc_hd__or2_1 _10112_ (.A(\sha256cu.msg_scheduler.mreg_3[19] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04300_));
 sky130_fd_sc_hd__o211a_1 _10113_ (.A1(\sha256cu.msg_scheduler.mreg_2[19] ),
    .A2(_04288_),
    .B1(_04300_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00543_));
 sky130_fd_sc_hd__buf_2 _10114_ (.A(_04166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04301_));
 sky130_fd_sc_hd__or2_1 _10115_ (.A(\sha256cu.msg_scheduler.mreg_3[20] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04302_));
 sky130_fd_sc_hd__o211a_1 _10116_ (.A1(\sha256cu.msg_scheduler.mreg_2[20] ),
    .A2(_04301_),
    .B1(_04302_),
    .C1(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00544_));
 sky130_fd_sc_hd__or2_1 _10117_ (.A(\sha256cu.msg_scheduler.mreg_3[21] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04303_));
 sky130_fd_sc_hd__buf_2 _10118_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04304_));
 sky130_fd_sc_hd__o211a_1 _10119_ (.A1(\sha256cu.msg_scheduler.mreg_2[21] ),
    .A2(_04301_),
    .B1(_04303_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00545_));
 sky130_fd_sc_hd__or2_1 _10120_ (.A(\sha256cu.msg_scheduler.mreg_3[22] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04305_));
 sky130_fd_sc_hd__o211a_1 _10121_ (.A1(\sha256cu.msg_scheduler.mreg_2[22] ),
    .A2(_04301_),
    .B1(_04305_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00546_));
 sky130_fd_sc_hd__or2_1 _10122_ (.A(\sha256cu.msg_scheduler.mreg_3[23] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04306_));
 sky130_fd_sc_hd__o211a_1 _10123_ (.A1(\sha256cu.msg_scheduler.mreg_2[23] ),
    .A2(_04301_),
    .B1(_04306_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _10124_ (.A(\sha256cu.msg_scheduler.mreg_3[24] ),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04307_));
 sky130_fd_sc_hd__o211a_1 _10125_ (.A1(\sha256cu.msg_scheduler.mreg_2[24] ),
    .A2(_04301_),
    .B1(_04307_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00548_));
 sky130_fd_sc_hd__clkbuf_2 _10126_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04308_));
 sky130_fd_sc_hd__or2_1 _10127_ (.A(\sha256cu.msg_scheduler.mreg_3[25] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04309_));
 sky130_fd_sc_hd__o211a_1 _10128_ (.A1(\sha256cu.msg_scheduler.mreg_2[25] ),
    .A2(_04301_),
    .B1(_04309_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00549_));
 sky130_fd_sc_hd__or2_1 _10129_ (.A(\sha256cu.msg_scheduler.mreg_3[26] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04310_));
 sky130_fd_sc_hd__o211a_1 _10130_ (.A1(\sha256cu.msg_scheduler.mreg_2[26] ),
    .A2(_04301_),
    .B1(_04310_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00550_));
 sky130_fd_sc_hd__or2_1 _10131_ (.A(\sha256cu.msg_scheduler.mreg_3[27] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04311_));
 sky130_fd_sc_hd__o211a_1 _10132_ (.A1(\sha256cu.msg_scheduler.mreg_2[27] ),
    .A2(_04301_),
    .B1(_04311_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00551_));
 sky130_fd_sc_hd__or2_1 _10133_ (.A(\sha256cu.msg_scheduler.mreg_3[28] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04312_));
 sky130_fd_sc_hd__o211a_1 _10134_ (.A1(\sha256cu.msg_scheduler.mreg_2[28] ),
    .A2(_04301_),
    .B1(_04312_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00552_));
 sky130_fd_sc_hd__or2_1 _10135_ (.A(\sha256cu.msg_scheduler.mreg_3[29] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04313_));
 sky130_fd_sc_hd__o211a_1 _10136_ (.A1(\sha256cu.msg_scheduler.mreg_2[29] ),
    .A2(_04301_),
    .B1(_04313_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00553_));
 sky130_fd_sc_hd__buf_2 _10137_ (.A(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04314_));
 sky130_fd_sc_hd__buf_2 _10138_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04315_));
 sky130_fd_sc_hd__or2_1 _10139_ (.A(\sha256cu.msg_scheduler.mreg_3[30] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04316_));
 sky130_fd_sc_hd__o211a_1 _10140_ (.A1(\sha256cu.msg_scheduler.mreg_2[30] ),
    .A2(_04315_),
    .B1(_04316_),
    .C1(_04304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _10141_ (.A(\sha256cu.msg_scheduler.mreg_3[31] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_4 _10142_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04318_));
 sky130_fd_sc_hd__o211a_1 _10143_ (.A1(\sha256cu.msg_scheduler.mreg_2[31] ),
    .A2(_04315_),
    .B1(_04317_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00555_));
 sky130_fd_sc_hd__or2_1 _10144_ (.A(\sha256cu.msg_scheduler.mreg_4[0] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04319_));
 sky130_fd_sc_hd__o211a_1 _10145_ (.A1(\sha256cu.msg_scheduler.mreg_3[0] ),
    .A2(_04315_),
    .B1(_04319_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00556_));
 sky130_fd_sc_hd__or2_1 _10146_ (.A(\sha256cu.msg_scheduler.mreg_4[1] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04320_));
 sky130_fd_sc_hd__o211a_1 _10147_ (.A1(\sha256cu.msg_scheduler.mreg_3[1] ),
    .A2(_04315_),
    .B1(_04320_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00557_));
 sky130_fd_sc_hd__or2_1 _10148_ (.A(\sha256cu.msg_scheduler.mreg_4[2] ),
    .B(_04308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04321_));
 sky130_fd_sc_hd__o211a_1 _10149_ (.A1(\sha256cu.msg_scheduler.mreg_3[2] ),
    .A2(_04315_),
    .B1(_04321_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00558_));
 sky130_fd_sc_hd__clkbuf_2 _10150_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04322_));
 sky130_fd_sc_hd__or2_1 _10151_ (.A(\sha256cu.msg_scheduler.mreg_4[3] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04323_));
 sky130_fd_sc_hd__o211a_1 _10152_ (.A1(\sha256cu.msg_scheduler.mreg_3[3] ),
    .A2(_04315_),
    .B1(_04323_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00559_));
 sky130_fd_sc_hd__or2_1 _10153_ (.A(\sha256cu.msg_scheduler.mreg_4[4] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04324_));
 sky130_fd_sc_hd__o211a_1 _10154_ (.A1(\sha256cu.msg_scheduler.mreg_3[4] ),
    .A2(_04315_),
    .B1(_04324_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _10155_ (.A(\sha256cu.msg_scheduler.mreg_4[5] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04325_));
 sky130_fd_sc_hd__o211a_1 _10156_ (.A1(\sha256cu.msg_scheduler.mreg_3[5] ),
    .A2(_04315_),
    .B1(_04325_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00561_));
 sky130_fd_sc_hd__or2_1 _10157_ (.A(\sha256cu.msg_scheduler.mreg_4[6] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04326_));
 sky130_fd_sc_hd__o211a_1 _10158_ (.A1(\sha256cu.msg_scheduler.mreg_3[6] ),
    .A2(_04315_),
    .B1(_04326_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00562_));
 sky130_fd_sc_hd__or2_1 _10159_ (.A(\sha256cu.msg_scheduler.mreg_4[7] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04327_));
 sky130_fd_sc_hd__o211a_1 _10160_ (.A1(\sha256cu.msg_scheduler.mreg_3[7] ),
    .A2(_04315_),
    .B1(_04327_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00563_));
 sky130_fd_sc_hd__buf_2 _10161_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04328_));
 sky130_fd_sc_hd__or2_1 _10162_ (.A(\sha256cu.msg_scheduler.mreg_4[8] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04329_));
 sky130_fd_sc_hd__o211a_1 _10163_ (.A1(\sha256cu.msg_scheduler.mreg_3[8] ),
    .A2(_04328_),
    .B1(_04329_),
    .C1(_04318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00564_));
 sky130_fd_sc_hd__or2_1 _10164_ (.A(\sha256cu.msg_scheduler.mreg_4[9] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04330_));
 sky130_fd_sc_hd__buf_2 _10165_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04331_));
 sky130_fd_sc_hd__o211a_1 _10166_ (.A1(\sha256cu.msg_scheduler.mreg_3[9] ),
    .A2(_04328_),
    .B1(_04330_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00565_));
 sky130_fd_sc_hd__or2_1 _10167_ (.A(\sha256cu.msg_scheduler.mreg_4[10] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04332_));
 sky130_fd_sc_hd__o211a_1 _10168_ (.A1(\sha256cu.msg_scheduler.mreg_3[10] ),
    .A2(_04328_),
    .B1(_04332_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00566_));
 sky130_fd_sc_hd__or2_1 _10169_ (.A(\sha256cu.msg_scheduler.mreg_4[11] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04333_));
 sky130_fd_sc_hd__o211a_1 _10170_ (.A1(\sha256cu.msg_scheduler.mreg_3[11] ),
    .A2(_04328_),
    .B1(_04333_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00567_));
 sky130_fd_sc_hd__or2_1 _10171_ (.A(\sha256cu.msg_scheduler.mreg_4[12] ),
    .B(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04334_));
 sky130_fd_sc_hd__o211a_1 _10172_ (.A1(\sha256cu.msg_scheduler.mreg_3[12] ),
    .A2(_04328_),
    .B1(_04334_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00568_));
 sky130_fd_sc_hd__clkbuf_2 _10173_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04335_));
 sky130_fd_sc_hd__or2_1 _10174_ (.A(\sha256cu.msg_scheduler.mreg_4[13] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04336_));
 sky130_fd_sc_hd__o211a_1 _10175_ (.A1(\sha256cu.msg_scheduler.mreg_3[13] ),
    .A2(_04328_),
    .B1(_04336_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00569_));
 sky130_fd_sc_hd__or2_1 _10176_ (.A(\sha256cu.msg_scheduler.mreg_4[14] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04337_));
 sky130_fd_sc_hd__o211a_1 _10177_ (.A1(\sha256cu.msg_scheduler.mreg_3[14] ),
    .A2(_04328_),
    .B1(_04337_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00570_));
 sky130_fd_sc_hd__or2_1 _10178_ (.A(\sha256cu.msg_scheduler.mreg_4[15] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04338_));
 sky130_fd_sc_hd__o211a_1 _10179_ (.A1(\sha256cu.msg_scheduler.mreg_3[15] ),
    .A2(_04328_),
    .B1(_04338_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00571_));
 sky130_fd_sc_hd__or2_1 _10180_ (.A(\sha256cu.msg_scheduler.mreg_4[16] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04339_));
 sky130_fd_sc_hd__o211a_1 _10181_ (.A1(\sha256cu.msg_scheduler.mreg_3[16] ),
    .A2(_04328_),
    .B1(_04339_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00572_));
 sky130_fd_sc_hd__or2_1 _10182_ (.A(\sha256cu.msg_scheduler.mreg_4[17] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04340_));
 sky130_fd_sc_hd__o211a_1 _10183_ (.A1(\sha256cu.msg_scheduler.mreg_3[17] ),
    .A2(_04328_),
    .B1(_04340_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00573_));
 sky130_fd_sc_hd__buf_2 _10184_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04341_));
 sky130_fd_sc_hd__or2_1 _10185_ (.A(\sha256cu.msg_scheduler.mreg_4[18] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04342_));
 sky130_fd_sc_hd__o211a_1 _10186_ (.A1(\sha256cu.msg_scheduler.mreg_3[18] ),
    .A2(_04341_),
    .B1(_04342_),
    .C1(_04331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00574_));
 sky130_fd_sc_hd__or2_1 _10187_ (.A(\sha256cu.msg_scheduler.mreg_4[19] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04343_));
 sky130_fd_sc_hd__buf_2 _10188_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04344_));
 sky130_fd_sc_hd__o211a_1 _10189_ (.A1(\sha256cu.msg_scheduler.mreg_3[19] ),
    .A2(_04341_),
    .B1(_04343_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00575_));
 sky130_fd_sc_hd__or2_1 _10190_ (.A(\sha256cu.msg_scheduler.mreg_4[20] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04345_));
 sky130_fd_sc_hd__o211a_1 _10191_ (.A1(\sha256cu.msg_scheduler.mreg_3[20] ),
    .A2(_04341_),
    .B1(_04345_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00576_));
 sky130_fd_sc_hd__or2_1 _10192_ (.A(\sha256cu.msg_scheduler.mreg_4[21] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04346_));
 sky130_fd_sc_hd__o211a_1 _10193_ (.A1(\sha256cu.msg_scheduler.mreg_3[21] ),
    .A2(_04341_),
    .B1(_04346_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00577_));
 sky130_fd_sc_hd__or2_1 _10194_ (.A(\sha256cu.msg_scheduler.mreg_4[22] ),
    .B(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04347_));
 sky130_fd_sc_hd__o211a_1 _10195_ (.A1(\sha256cu.msg_scheduler.mreg_3[22] ),
    .A2(_04341_),
    .B1(_04347_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00578_));
 sky130_fd_sc_hd__clkbuf_2 _10196_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04348_));
 sky130_fd_sc_hd__or2_1 _10197_ (.A(\sha256cu.msg_scheduler.mreg_4[23] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04349_));
 sky130_fd_sc_hd__o211a_1 _10198_ (.A1(\sha256cu.msg_scheduler.mreg_3[23] ),
    .A2(_04341_),
    .B1(_04349_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00579_));
 sky130_fd_sc_hd__or2_1 _10199_ (.A(\sha256cu.msg_scheduler.mreg_4[24] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04350_));
 sky130_fd_sc_hd__o211a_1 _10200_ (.A1(\sha256cu.msg_scheduler.mreg_3[24] ),
    .A2(_04341_),
    .B1(_04350_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00580_));
 sky130_fd_sc_hd__or2_1 _10201_ (.A(\sha256cu.msg_scheduler.mreg_4[25] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04351_));
 sky130_fd_sc_hd__o211a_1 _10202_ (.A1(\sha256cu.msg_scheduler.mreg_3[25] ),
    .A2(_04341_),
    .B1(_04351_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00581_));
 sky130_fd_sc_hd__or2_1 _10203_ (.A(\sha256cu.msg_scheduler.mreg_4[26] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04352_));
 sky130_fd_sc_hd__o211a_1 _10204_ (.A1(\sha256cu.msg_scheduler.mreg_3[26] ),
    .A2(_04341_),
    .B1(_04352_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00582_));
 sky130_fd_sc_hd__or2_1 _10205_ (.A(\sha256cu.msg_scheduler.mreg_4[27] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04353_));
 sky130_fd_sc_hd__o211a_1 _10206_ (.A1(\sha256cu.msg_scheduler.mreg_3[27] ),
    .A2(_04341_),
    .B1(_04353_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00583_));
 sky130_fd_sc_hd__buf_2 _10207_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04354_));
 sky130_fd_sc_hd__or2_1 _10208_ (.A(\sha256cu.msg_scheduler.mreg_4[28] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04355_));
 sky130_fd_sc_hd__o211a_1 _10209_ (.A1(\sha256cu.msg_scheduler.mreg_3[28] ),
    .A2(_04354_),
    .B1(_04355_),
    .C1(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00584_));
 sky130_fd_sc_hd__or2_1 _10210_ (.A(\sha256cu.msg_scheduler.mreg_4[29] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04356_));
 sky130_fd_sc_hd__buf_2 _10211_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04357_));
 sky130_fd_sc_hd__o211a_1 _10212_ (.A1(\sha256cu.msg_scheduler.mreg_3[29] ),
    .A2(_04354_),
    .B1(_04356_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00585_));
 sky130_fd_sc_hd__or2_1 _10213_ (.A(\sha256cu.msg_scheduler.mreg_4[30] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04358_));
 sky130_fd_sc_hd__o211a_1 _10214_ (.A1(\sha256cu.msg_scheduler.mreg_3[30] ),
    .A2(_04354_),
    .B1(_04358_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00586_));
 sky130_fd_sc_hd__or2_1 _10215_ (.A(\sha256cu.msg_scheduler.mreg_4[31] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04359_));
 sky130_fd_sc_hd__o211a_1 _10216_ (.A1(\sha256cu.msg_scheduler.mreg_3[31] ),
    .A2(_04354_),
    .B1(_04359_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00587_));
 sky130_fd_sc_hd__or2_1 _10217_ (.A(\sha256cu.msg_scheduler.mreg_5[0] ),
    .B(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04360_));
 sky130_fd_sc_hd__o211a_1 _10218_ (.A1(\sha256cu.msg_scheduler.mreg_4[0] ),
    .A2(_04354_),
    .B1(_04360_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00588_));
 sky130_fd_sc_hd__clkbuf_2 _10219_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04361_));
 sky130_fd_sc_hd__or2_1 _10220_ (.A(\sha256cu.msg_scheduler.mreg_5[1] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04362_));
 sky130_fd_sc_hd__o211a_1 _10221_ (.A1(\sha256cu.msg_scheduler.mreg_4[1] ),
    .A2(_04354_),
    .B1(_04362_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00589_));
 sky130_fd_sc_hd__or2_1 _10222_ (.A(\sha256cu.msg_scheduler.mreg_5[2] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04363_));
 sky130_fd_sc_hd__o211a_1 _10223_ (.A1(\sha256cu.msg_scheduler.mreg_4[2] ),
    .A2(_04354_),
    .B1(_04363_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00590_));
 sky130_fd_sc_hd__or2_1 _10224_ (.A(\sha256cu.msg_scheduler.mreg_5[3] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04364_));
 sky130_fd_sc_hd__o211a_1 _10225_ (.A1(\sha256cu.msg_scheduler.mreg_4[3] ),
    .A2(_04354_),
    .B1(_04364_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00591_));
 sky130_fd_sc_hd__or2_1 _10226_ (.A(\sha256cu.msg_scheduler.mreg_5[4] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04365_));
 sky130_fd_sc_hd__o211a_1 _10227_ (.A1(\sha256cu.msg_scheduler.mreg_4[4] ),
    .A2(_04354_),
    .B1(_04365_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00592_));
 sky130_fd_sc_hd__or2_1 _10228_ (.A(\sha256cu.msg_scheduler.mreg_5[5] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04366_));
 sky130_fd_sc_hd__o211a_1 _10229_ (.A1(\sha256cu.msg_scheduler.mreg_4[5] ),
    .A2(_04354_),
    .B1(_04366_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00593_));
 sky130_fd_sc_hd__buf_2 _10230_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04367_));
 sky130_fd_sc_hd__or2_1 _10231_ (.A(\sha256cu.msg_scheduler.mreg_5[6] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04368_));
 sky130_fd_sc_hd__o211a_1 _10232_ (.A1(\sha256cu.msg_scheduler.mreg_4[6] ),
    .A2(_04367_),
    .B1(_04368_),
    .C1(_04357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00594_));
 sky130_fd_sc_hd__or2_1 _10233_ (.A(\sha256cu.msg_scheduler.mreg_5[7] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04369_));
 sky130_fd_sc_hd__buf_2 _10234_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04370_));
 sky130_fd_sc_hd__o211a_1 _10235_ (.A1(\sha256cu.msg_scheduler.mreg_4[7] ),
    .A2(_04367_),
    .B1(_04369_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00595_));
 sky130_fd_sc_hd__or2_1 _10236_ (.A(\sha256cu.msg_scheduler.mreg_5[8] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04371_));
 sky130_fd_sc_hd__o211a_1 _10237_ (.A1(\sha256cu.msg_scheduler.mreg_4[8] ),
    .A2(_04367_),
    .B1(_04371_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00596_));
 sky130_fd_sc_hd__or2_1 _10238_ (.A(\sha256cu.msg_scheduler.mreg_5[9] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04372_));
 sky130_fd_sc_hd__o211a_1 _10239_ (.A1(\sha256cu.msg_scheduler.mreg_4[9] ),
    .A2(_04367_),
    .B1(_04372_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00597_));
 sky130_fd_sc_hd__or2_1 _10240_ (.A(\sha256cu.msg_scheduler.mreg_5[10] ),
    .B(_04361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04373_));
 sky130_fd_sc_hd__o211a_1 _10241_ (.A1(\sha256cu.msg_scheduler.mreg_4[10] ),
    .A2(_04367_),
    .B1(_04373_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00598_));
 sky130_fd_sc_hd__clkbuf_2 _10242_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04374_));
 sky130_fd_sc_hd__or2_1 _10243_ (.A(\sha256cu.msg_scheduler.mreg_5[11] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04375_));
 sky130_fd_sc_hd__o211a_1 _10244_ (.A1(\sha256cu.msg_scheduler.mreg_4[11] ),
    .A2(_04367_),
    .B1(_04375_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00599_));
 sky130_fd_sc_hd__or2_1 _10245_ (.A(\sha256cu.msg_scheduler.mreg_5[12] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04376_));
 sky130_fd_sc_hd__o211a_1 _10246_ (.A1(\sha256cu.msg_scheduler.mreg_4[12] ),
    .A2(_04367_),
    .B1(_04376_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00600_));
 sky130_fd_sc_hd__or2_1 _10247_ (.A(\sha256cu.msg_scheduler.mreg_5[13] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04377_));
 sky130_fd_sc_hd__o211a_1 _10248_ (.A1(\sha256cu.msg_scheduler.mreg_4[13] ),
    .A2(_04367_),
    .B1(_04377_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00601_));
 sky130_fd_sc_hd__or2_1 _10249_ (.A(\sha256cu.msg_scheduler.mreg_5[14] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04378_));
 sky130_fd_sc_hd__o211a_1 _10250_ (.A1(\sha256cu.msg_scheduler.mreg_4[14] ),
    .A2(_04367_),
    .B1(_04378_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00602_));
 sky130_fd_sc_hd__or2_1 _10251_ (.A(\sha256cu.msg_scheduler.mreg_5[15] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04379_));
 sky130_fd_sc_hd__o211a_1 _10252_ (.A1(\sha256cu.msg_scheduler.mreg_4[15] ),
    .A2(_04367_),
    .B1(_04379_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00603_));
 sky130_fd_sc_hd__buf_2 _10253_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04380_));
 sky130_fd_sc_hd__or2_1 _10254_ (.A(\sha256cu.msg_scheduler.mreg_5[16] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04381_));
 sky130_fd_sc_hd__o211a_1 _10255_ (.A1(\sha256cu.msg_scheduler.mreg_4[16] ),
    .A2(_04380_),
    .B1(_04381_),
    .C1(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00604_));
 sky130_fd_sc_hd__or2_1 _10256_ (.A(\sha256cu.msg_scheduler.mreg_5[17] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04382_));
 sky130_fd_sc_hd__buf_2 _10257_ (.A(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04383_));
 sky130_fd_sc_hd__o211a_1 _10258_ (.A1(\sha256cu.msg_scheduler.mreg_4[17] ),
    .A2(_04380_),
    .B1(_04382_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00605_));
 sky130_fd_sc_hd__or2_1 _10259_ (.A(\sha256cu.msg_scheduler.mreg_5[18] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04384_));
 sky130_fd_sc_hd__o211a_1 _10260_ (.A1(\sha256cu.msg_scheduler.mreg_4[18] ),
    .A2(_04380_),
    .B1(_04384_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00606_));
 sky130_fd_sc_hd__or2_1 _10261_ (.A(\sha256cu.msg_scheduler.mreg_5[19] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04385_));
 sky130_fd_sc_hd__o211a_1 _10262_ (.A1(\sha256cu.msg_scheduler.mreg_4[19] ),
    .A2(_04380_),
    .B1(_04385_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00607_));
 sky130_fd_sc_hd__or2_1 _10263_ (.A(\sha256cu.msg_scheduler.mreg_5[20] ),
    .B(_04374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04386_));
 sky130_fd_sc_hd__o211a_1 _10264_ (.A1(\sha256cu.msg_scheduler.mreg_4[20] ),
    .A2(_04380_),
    .B1(_04386_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00608_));
 sky130_fd_sc_hd__clkbuf_2 _10265_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04387_));
 sky130_fd_sc_hd__or2_1 _10266_ (.A(\sha256cu.msg_scheduler.mreg_5[21] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04388_));
 sky130_fd_sc_hd__o211a_1 _10267_ (.A1(\sha256cu.msg_scheduler.mreg_4[21] ),
    .A2(_04380_),
    .B1(_04388_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00609_));
 sky130_fd_sc_hd__or2_1 _10268_ (.A(\sha256cu.msg_scheduler.mreg_5[22] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04389_));
 sky130_fd_sc_hd__o211a_1 _10269_ (.A1(\sha256cu.msg_scheduler.mreg_4[22] ),
    .A2(_04380_),
    .B1(_04389_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00610_));
 sky130_fd_sc_hd__or2_1 _10270_ (.A(\sha256cu.msg_scheduler.mreg_5[23] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04390_));
 sky130_fd_sc_hd__o211a_1 _10271_ (.A1(\sha256cu.msg_scheduler.mreg_4[23] ),
    .A2(_04380_),
    .B1(_04390_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00611_));
 sky130_fd_sc_hd__or2_1 _10272_ (.A(\sha256cu.msg_scheduler.mreg_5[24] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04391_));
 sky130_fd_sc_hd__o211a_1 _10273_ (.A1(\sha256cu.msg_scheduler.mreg_4[24] ),
    .A2(_04380_),
    .B1(_04391_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00612_));
 sky130_fd_sc_hd__or2_1 _10274_ (.A(\sha256cu.msg_scheduler.mreg_5[25] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04392_));
 sky130_fd_sc_hd__o211a_1 _10275_ (.A1(\sha256cu.msg_scheduler.mreg_4[25] ),
    .A2(_04380_),
    .B1(_04392_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00613_));
 sky130_fd_sc_hd__buf_2 _10276_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04393_));
 sky130_fd_sc_hd__or2_1 _10277_ (.A(\sha256cu.msg_scheduler.mreg_5[26] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04394_));
 sky130_fd_sc_hd__o211a_1 _10278_ (.A1(\sha256cu.msg_scheduler.mreg_4[26] ),
    .A2(_04393_),
    .B1(_04394_),
    .C1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00614_));
 sky130_fd_sc_hd__or2_1 _10279_ (.A(\sha256cu.msg_scheduler.mreg_5[27] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04395_));
 sky130_fd_sc_hd__buf_2 _10280_ (.A(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04396_));
 sky130_fd_sc_hd__buf_2 _10281_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04397_));
 sky130_fd_sc_hd__o211a_1 _10282_ (.A1(\sha256cu.msg_scheduler.mreg_4[27] ),
    .A2(_04393_),
    .B1(_04395_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00615_));
 sky130_fd_sc_hd__or2_1 _10283_ (.A(\sha256cu.msg_scheduler.mreg_5[28] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04398_));
 sky130_fd_sc_hd__o211a_1 _10284_ (.A1(\sha256cu.msg_scheduler.mreg_4[28] ),
    .A2(_04393_),
    .B1(_04398_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00616_));
 sky130_fd_sc_hd__or2_1 _10285_ (.A(\sha256cu.msg_scheduler.mreg_5[29] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04399_));
 sky130_fd_sc_hd__o211a_1 _10286_ (.A1(\sha256cu.msg_scheduler.mreg_4[29] ),
    .A2(_04393_),
    .B1(_04399_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00617_));
 sky130_fd_sc_hd__or2_1 _10287_ (.A(\sha256cu.msg_scheduler.mreg_5[30] ),
    .B(_04387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04400_));
 sky130_fd_sc_hd__o211a_1 _10288_ (.A1(\sha256cu.msg_scheduler.mreg_4[30] ),
    .A2(_04393_),
    .B1(_04400_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00618_));
 sky130_fd_sc_hd__clkbuf_2 _10289_ (.A(_04281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04401_));
 sky130_fd_sc_hd__or2_1 _10290_ (.A(\sha256cu.msg_scheduler.mreg_5[31] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04402_));
 sky130_fd_sc_hd__o211a_1 _10291_ (.A1(\sha256cu.msg_scheduler.mreg_4[31] ),
    .A2(_04393_),
    .B1(_04402_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00619_));
 sky130_fd_sc_hd__or2_1 _10292_ (.A(\sha256cu.msg_scheduler.mreg_6[0] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04403_));
 sky130_fd_sc_hd__o211a_1 _10293_ (.A1(\sha256cu.msg_scheduler.mreg_5[0] ),
    .A2(_04393_),
    .B1(_04403_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00620_));
 sky130_fd_sc_hd__or2_1 _10294_ (.A(\sha256cu.msg_scheduler.mreg_6[1] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04404_));
 sky130_fd_sc_hd__o211a_1 _10295_ (.A1(\sha256cu.msg_scheduler.mreg_5[1] ),
    .A2(_04393_),
    .B1(_04404_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00621_));
 sky130_fd_sc_hd__or2_1 _10296_ (.A(\sha256cu.msg_scheduler.mreg_6[2] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04405_));
 sky130_fd_sc_hd__o211a_1 _10297_ (.A1(\sha256cu.msg_scheduler.mreg_5[2] ),
    .A2(_04393_),
    .B1(_04405_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00622_));
 sky130_fd_sc_hd__or2_1 _10298_ (.A(\sha256cu.msg_scheduler.mreg_6[3] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04406_));
 sky130_fd_sc_hd__o211a_1 _10299_ (.A1(\sha256cu.msg_scheduler.mreg_5[3] ),
    .A2(_04393_),
    .B1(_04406_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00623_));
 sky130_fd_sc_hd__buf_2 _10300_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04407_));
 sky130_fd_sc_hd__or2_1 _10301_ (.A(\sha256cu.msg_scheduler.mreg_6[4] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04408_));
 sky130_fd_sc_hd__o211a_1 _10302_ (.A1(\sha256cu.msg_scheduler.mreg_5[4] ),
    .A2(_04407_),
    .B1(_04408_),
    .C1(_04397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00624_));
 sky130_fd_sc_hd__or2_1 _10303_ (.A(\sha256cu.msg_scheduler.mreg_6[5] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04409_));
 sky130_fd_sc_hd__buf_2 _10304_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04410_));
 sky130_fd_sc_hd__o211a_1 _10305_ (.A1(\sha256cu.msg_scheduler.mreg_5[5] ),
    .A2(_04407_),
    .B1(_04409_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00625_));
 sky130_fd_sc_hd__or2_1 _10306_ (.A(\sha256cu.msg_scheduler.mreg_6[6] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04411_));
 sky130_fd_sc_hd__o211a_1 _10307_ (.A1(\sha256cu.msg_scheduler.mreg_5[6] ),
    .A2(_04407_),
    .B1(_04411_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00626_));
 sky130_fd_sc_hd__or2_1 _10308_ (.A(\sha256cu.msg_scheduler.mreg_6[7] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04412_));
 sky130_fd_sc_hd__o211a_1 _10309_ (.A1(\sha256cu.msg_scheduler.mreg_5[7] ),
    .A2(_04407_),
    .B1(_04412_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00627_));
 sky130_fd_sc_hd__or2_1 _10310_ (.A(\sha256cu.msg_scheduler.mreg_6[8] ),
    .B(_04401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04413_));
 sky130_fd_sc_hd__o211a_1 _10311_ (.A1(\sha256cu.msg_scheduler.mreg_5[8] ),
    .A2(_04407_),
    .B1(_04413_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00628_));
 sky130_fd_sc_hd__clkbuf_4 _10312_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_2 _10313_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04415_));
 sky130_fd_sc_hd__or2_1 _10314_ (.A(\sha256cu.msg_scheduler.mreg_6[9] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04416_));
 sky130_fd_sc_hd__o211a_1 _10315_ (.A1(\sha256cu.msg_scheduler.mreg_5[9] ),
    .A2(_04407_),
    .B1(_04416_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00629_));
 sky130_fd_sc_hd__or2_1 _10316_ (.A(\sha256cu.msg_scheduler.mreg_6[10] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04417_));
 sky130_fd_sc_hd__o211a_1 _10317_ (.A1(\sha256cu.msg_scheduler.mreg_5[10] ),
    .A2(_04407_),
    .B1(_04417_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00630_));
 sky130_fd_sc_hd__or2_1 _10318_ (.A(\sha256cu.msg_scheduler.mreg_6[11] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04418_));
 sky130_fd_sc_hd__o211a_1 _10319_ (.A1(\sha256cu.msg_scheduler.mreg_5[11] ),
    .A2(_04407_),
    .B1(_04418_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00631_));
 sky130_fd_sc_hd__or2_1 _10320_ (.A(\sha256cu.msg_scheduler.mreg_6[12] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04419_));
 sky130_fd_sc_hd__o211a_1 _10321_ (.A1(\sha256cu.msg_scheduler.mreg_5[12] ),
    .A2(_04407_),
    .B1(_04419_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00632_));
 sky130_fd_sc_hd__or2_1 _10322_ (.A(\sha256cu.msg_scheduler.mreg_6[13] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04420_));
 sky130_fd_sc_hd__o211a_1 _10323_ (.A1(\sha256cu.msg_scheduler.mreg_5[13] ),
    .A2(_04407_),
    .B1(_04420_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00633_));
 sky130_fd_sc_hd__buf_2 _10324_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04421_));
 sky130_fd_sc_hd__or2_1 _10325_ (.A(\sha256cu.msg_scheduler.mreg_6[14] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04422_));
 sky130_fd_sc_hd__o211a_1 _10326_ (.A1(\sha256cu.msg_scheduler.mreg_5[14] ),
    .A2(_04421_),
    .B1(_04422_),
    .C1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00634_));
 sky130_fd_sc_hd__or2_1 _10327_ (.A(\sha256cu.msg_scheduler.mreg_6[15] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04423_));
 sky130_fd_sc_hd__buf_2 _10328_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04424_));
 sky130_fd_sc_hd__o211a_1 _10329_ (.A1(\sha256cu.msg_scheduler.mreg_5[15] ),
    .A2(_04421_),
    .B1(_04423_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00635_));
 sky130_fd_sc_hd__or2_1 _10330_ (.A(\sha256cu.msg_scheduler.mreg_6[16] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04425_));
 sky130_fd_sc_hd__o211a_1 _10331_ (.A1(\sha256cu.msg_scheduler.mreg_5[16] ),
    .A2(_04421_),
    .B1(_04425_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00636_));
 sky130_fd_sc_hd__or2_1 _10332_ (.A(\sha256cu.msg_scheduler.mreg_6[17] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04426_));
 sky130_fd_sc_hd__o211a_1 _10333_ (.A1(\sha256cu.msg_scheduler.mreg_5[17] ),
    .A2(_04421_),
    .B1(_04426_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00637_));
 sky130_fd_sc_hd__or2_1 _10334_ (.A(\sha256cu.msg_scheduler.mreg_6[18] ),
    .B(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04427_));
 sky130_fd_sc_hd__o211a_1 _10335_ (.A1(\sha256cu.msg_scheduler.mreg_5[18] ),
    .A2(_04421_),
    .B1(_04427_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00638_));
 sky130_fd_sc_hd__clkbuf_2 _10336_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04428_));
 sky130_fd_sc_hd__or2_1 _10337_ (.A(\sha256cu.msg_scheduler.mreg_6[19] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04429_));
 sky130_fd_sc_hd__o211a_1 _10338_ (.A1(\sha256cu.msg_scheduler.mreg_5[19] ),
    .A2(_04421_),
    .B1(_04429_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00639_));
 sky130_fd_sc_hd__or2_1 _10339_ (.A(\sha256cu.msg_scheduler.mreg_6[20] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04430_));
 sky130_fd_sc_hd__o211a_1 _10340_ (.A1(\sha256cu.msg_scheduler.mreg_5[20] ),
    .A2(_04421_),
    .B1(_04430_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00640_));
 sky130_fd_sc_hd__or2_1 _10341_ (.A(\sha256cu.msg_scheduler.mreg_6[21] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04431_));
 sky130_fd_sc_hd__o211a_1 _10342_ (.A1(\sha256cu.msg_scheduler.mreg_5[21] ),
    .A2(_04421_),
    .B1(_04431_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00641_));
 sky130_fd_sc_hd__or2_1 _10343_ (.A(\sha256cu.msg_scheduler.mreg_6[22] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04432_));
 sky130_fd_sc_hd__o211a_1 _10344_ (.A1(\sha256cu.msg_scheduler.mreg_5[22] ),
    .A2(_04421_),
    .B1(_04432_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00642_));
 sky130_fd_sc_hd__or2_1 _10345_ (.A(\sha256cu.msg_scheduler.mreg_6[23] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04433_));
 sky130_fd_sc_hd__o211a_1 _10346_ (.A1(\sha256cu.msg_scheduler.mreg_5[23] ),
    .A2(_04421_),
    .B1(_04433_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00643_));
 sky130_fd_sc_hd__clkbuf_4 _10347_ (.A(_04314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04434_));
 sky130_fd_sc_hd__or2_1 _10348_ (.A(\sha256cu.msg_scheduler.mreg_6[24] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04435_));
 sky130_fd_sc_hd__o211a_1 _10349_ (.A1(\sha256cu.msg_scheduler.mreg_5[24] ),
    .A2(_04434_),
    .B1(_04435_),
    .C1(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00644_));
 sky130_fd_sc_hd__or2_1 _10350_ (.A(\sha256cu.msg_scheduler.mreg_6[25] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04436_));
 sky130_fd_sc_hd__buf_2 _10351_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04437_));
 sky130_fd_sc_hd__o211a_1 _10352_ (.A1(\sha256cu.msg_scheduler.mreg_5[25] ),
    .A2(_04434_),
    .B1(_04436_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00645_));
 sky130_fd_sc_hd__or2_1 _10353_ (.A(\sha256cu.msg_scheduler.mreg_6[26] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04438_));
 sky130_fd_sc_hd__o211a_1 _10354_ (.A1(\sha256cu.msg_scheduler.mreg_5[26] ),
    .A2(_04434_),
    .B1(_04438_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00646_));
 sky130_fd_sc_hd__or2_1 _10355_ (.A(\sha256cu.msg_scheduler.mreg_6[27] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04439_));
 sky130_fd_sc_hd__o211a_1 _10356_ (.A1(\sha256cu.msg_scheduler.mreg_5[27] ),
    .A2(_04434_),
    .B1(_04439_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00647_));
 sky130_fd_sc_hd__or2_1 _10357_ (.A(\sha256cu.msg_scheduler.mreg_6[28] ),
    .B(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04440_));
 sky130_fd_sc_hd__o211a_1 _10358_ (.A1(\sha256cu.msg_scheduler.mreg_5[28] ),
    .A2(_04434_),
    .B1(_04440_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00648_));
 sky130_fd_sc_hd__clkbuf_2 _10359_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04441_));
 sky130_fd_sc_hd__or2_1 _10360_ (.A(\sha256cu.msg_scheduler.mreg_6[29] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04442_));
 sky130_fd_sc_hd__o211a_1 _10361_ (.A1(\sha256cu.msg_scheduler.mreg_5[29] ),
    .A2(_04434_),
    .B1(_04442_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00649_));
 sky130_fd_sc_hd__or2_1 _10362_ (.A(\sha256cu.msg_scheduler.mreg_6[30] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04443_));
 sky130_fd_sc_hd__o211a_1 _10363_ (.A1(\sha256cu.msg_scheduler.mreg_5[30] ),
    .A2(_04434_),
    .B1(_04443_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00650_));
 sky130_fd_sc_hd__or2_1 _10364_ (.A(\sha256cu.msg_scheduler.mreg_6[31] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04444_));
 sky130_fd_sc_hd__o211a_1 _10365_ (.A1(\sha256cu.msg_scheduler.mreg_5[31] ),
    .A2(_04434_),
    .B1(_04444_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00651_));
 sky130_fd_sc_hd__or2_1 _10366_ (.A(\sha256cu.msg_scheduler.mreg_7[0] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04445_));
 sky130_fd_sc_hd__o211a_1 _10367_ (.A1(\sha256cu.msg_scheduler.mreg_6[0] ),
    .A2(_04434_),
    .B1(_04445_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00652_));
 sky130_fd_sc_hd__or2_1 _10368_ (.A(\sha256cu.msg_scheduler.mreg_7[1] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04446_));
 sky130_fd_sc_hd__o211a_1 _10369_ (.A1(\sha256cu.msg_scheduler.mreg_6[1] ),
    .A2(_04434_),
    .B1(_04446_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00653_));
 sky130_fd_sc_hd__clkbuf_4 _10370_ (.A(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04447_));
 sky130_fd_sc_hd__buf_2 _10371_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04448_));
 sky130_fd_sc_hd__or2_1 _10372_ (.A(\sha256cu.msg_scheduler.mreg_7[2] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04449_));
 sky130_fd_sc_hd__o211a_1 _10373_ (.A1(\sha256cu.msg_scheduler.mreg_6[2] ),
    .A2(_04448_),
    .B1(_04449_),
    .C1(_04437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00654_));
 sky130_fd_sc_hd__or2_1 _10374_ (.A(\sha256cu.msg_scheduler.mreg_7[3] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04450_));
 sky130_fd_sc_hd__buf_2 _10375_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04451_));
 sky130_fd_sc_hd__o211a_1 _10376_ (.A1(\sha256cu.msg_scheduler.mreg_6[3] ),
    .A2(_04448_),
    .B1(_04450_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00655_));
 sky130_fd_sc_hd__or2_1 _10377_ (.A(\sha256cu.msg_scheduler.mreg_7[4] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04452_));
 sky130_fd_sc_hd__o211a_1 _10378_ (.A1(\sha256cu.msg_scheduler.mreg_6[4] ),
    .A2(_04448_),
    .B1(_04452_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00656_));
 sky130_fd_sc_hd__or2_1 _10379_ (.A(\sha256cu.msg_scheduler.mreg_7[5] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04453_));
 sky130_fd_sc_hd__o211a_1 _10380_ (.A1(\sha256cu.msg_scheduler.mreg_6[5] ),
    .A2(_04448_),
    .B1(_04453_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00657_));
 sky130_fd_sc_hd__or2_1 _10381_ (.A(\sha256cu.msg_scheduler.mreg_7[6] ),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04454_));
 sky130_fd_sc_hd__o211a_1 _10382_ (.A1(\sha256cu.msg_scheduler.mreg_6[6] ),
    .A2(_04448_),
    .B1(_04454_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00658_));
 sky130_fd_sc_hd__clkbuf_2 _10383_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04455_));
 sky130_fd_sc_hd__or2_1 _10384_ (.A(\sha256cu.msg_scheduler.mreg_7[7] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04456_));
 sky130_fd_sc_hd__o211a_1 _10385_ (.A1(\sha256cu.msg_scheduler.mreg_6[7] ),
    .A2(_04448_),
    .B1(_04456_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00659_));
 sky130_fd_sc_hd__or2_1 _10386_ (.A(\sha256cu.msg_scheduler.mreg_7[8] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04457_));
 sky130_fd_sc_hd__o211a_1 _10387_ (.A1(\sha256cu.msg_scheduler.mreg_6[8] ),
    .A2(_04448_),
    .B1(_04457_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00660_));
 sky130_fd_sc_hd__or2_1 _10388_ (.A(\sha256cu.msg_scheduler.mreg_7[9] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04458_));
 sky130_fd_sc_hd__o211a_1 _10389_ (.A1(\sha256cu.msg_scheduler.mreg_6[9] ),
    .A2(_04448_),
    .B1(_04458_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00661_));
 sky130_fd_sc_hd__or2_1 _10390_ (.A(\sha256cu.msg_scheduler.mreg_7[10] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04459_));
 sky130_fd_sc_hd__o211a_1 _10391_ (.A1(\sha256cu.msg_scheduler.mreg_6[10] ),
    .A2(_04448_),
    .B1(_04459_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00662_));
 sky130_fd_sc_hd__or2_1 _10392_ (.A(\sha256cu.msg_scheduler.mreg_7[11] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04460_));
 sky130_fd_sc_hd__o211a_1 _10393_ (.A1(\sha256cu.msg_scheduler.mreg_6[11] ),
    .A2(_04448_),
    .B1(_04460_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00663_));
 sky130_fd_sc_hd__buf_2 _10394_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04461_));
 sky130_fd_sc_hd__or2_1 _10395_ (.A(\sha256cu.msg_scheduler.mreg_7[12] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04462_));
 sky130_fd_sc_hd__o211a_1 _10396_ (.A1(\sha256cu.msg_scheduler.mreg_6[12] ),
    .A2(_04461_),
    .B1(_04462_),
    .C1(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00664_));
 sky130_fd_sc_hd__or2_1 _10397_ (.A(\sha256cu.msg_scheduler.mreg_7[13] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04463_));
 sky130_fd_sc_hd__buf_2 _10398_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04464_));
 sky130_fd_sc_hd__o211a_1 _10399_ (.A1(\sha256cu.msg_scheduler.mreg_6[13] ),
    .A2(_04461_),
    .B1(_04463_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00665_));
 sky130_fd_sc_hd__or2_1 _10400_ (.A(\sha256cu.msg_scheduler.mreg_7[14] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04465_));
 sky130_fd_sc_hd__o211a_1 _10401_ (.A1(\sha256cu.msg_scheduler.mreg_6[14] ),
    .A2(_04461_),
    .B1(_04465_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00666_));
 sky130_fd_sc_hd__or2_1 _10402_ (.A(\sha256cu.msg_scheduler.mreg_7[15] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04466_));
 sky130_fd_sc_hd__o211a_1 _10403_ (.A1(\sha256cu.msg_scheduler.mreg_6[15] ),
    .A2(_04461_),
    .B1(_04466_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00667_));
 sky130_fd_sc_hd__or2_1 _10404_ (.A(\sha256cu.msg_scheduler.mreg_7[16] ),
    .B(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04467_));
 sky130_fd_sc_hd__o211a_1 _10405_ (.A1(\sha256cu.msg_scheduler.mreg_6[16] ),
    .A2(_04461_),
    .B1(_04467_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00668_));
 sky130_fd_sc_hd__clkbuf_2 _10406_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04468_));
 sky130_fd_sc_hd__or2_1 _10407_ (.A(\sha256cu.msg_scheduler.mreg_7[17] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04469_));
 sky130_fd_sc_hd__o211a_1 _10408_ (.A1(\sha256cu.msg_scheduler.mreg_6[17] ),
    .A2(_04461_),
    .B1(_04469_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00669_));
 sky130_fd_sc_hd__or2_1 _10409_ (.A(\sha256cu.msg_scheduler.mreg_7[18] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04470_));
 sky130_fd_sc_hd__o211a_1 _10410_ (.A1(\sha256cu.msg_scheduler.mreg_6[18] ),
    .A2(_04461_),
    .B1(_04470_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00670_));
 sky130_fd_sc_hd__or2_1 _10411_ (.A(\sha256cu.msg_scheduler.mreg_7[19] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04471_));
 sky130_fd_sc_hd__o211a_1 _10412_ (.A1(\sha256cu.msg_scheduler.mreg_6[19] ),
    .A2(_04461_),
    .B1(_04471_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00671_));
 sky130_fd_sc_hd__or2_1 _10413_ (.A(\sha256cu.msg_scheduler.mreg_7[20] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04472_));
 sky130_fd_sc_hd__o211a_1 _10414_ (.A1(\sha256cu.msg_scheduler.mreg_6[20] ),
    .A2(_04461_),
    .B1(_04472_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00672_));
 sky130_fd_sc_hd__or2_1 _10415_ (.A(\sha256cu.msg_scheduler.mreg_7[21] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04473_));
 sky130_fd_sc_hd__o211a_1 _10416_ (.A1(\sha256cu.msg_scheduler.mreg_6[21] ),
    .A2(_04461_),
    .B1(_04473_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00673_));
 sky130_fd_sc_hd__buf_2 _10417_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04474_));
 sky130_fd_sc_hd__or2_1 _10418_ (.A(\sha256cu.msg_scheduler.mreg_7[22] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04475_));
 sky130_fd_sc_hd__o211a_1 _10419_ (.A1(\sha256cu.msg_scheduler.mreg_6[22] ),
    .A2(_04474_),
    .B1(_04475_),
    .C1(_04464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00674_));
 sky130_fd_sc_hd__or2_1 _10420_ (.A(\sha256cu.msg_scheduler.mreg_7[23] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04476_));
 sky130_fd_sc_hd__buf_2 _10421_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04477_));
 sky130_fd_sc_hd__o211a_1 _10422_ (.A1(\sha256cu.msg_scheduler.mreg_6[23] ),
    .A2(_04474_),
    .B1(_04476_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00675_));
 sky130_fd_sc_hd__or2_1 _10423_ (.A(\sha256cu.msg_scheduler.mreg_7[24] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04478_));
 sky130_fd_sc_hd__o211a_1 _10424_ (.A1(\sha256cu.msg_scheduler.mreg_6[24] ),
    .A2(_04474_),
    .B1(_04478_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00676_));
 sky130_fd_sc_hd__or2_1 _10425_ (.A(\sha256cu.msg_scheduler.mreg_7[25] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04479_));
 sky130_fd_sc_hd__o211a_1 _10426_ (.A1(\sha256cu.msg_scheduler.mreg_6[25] ),
    .A2(_04474_),
    .B1(_04479_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00677_));
 sky130_fd_sc_hd__or2_1 _10427_ (.A(\sha256cu.msg_scheduler.mreg_7[26] ),
    .B(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04480_));
 sky130_fd_sc_hd__o211a_1 _10428_ (.A1(\sha256cu.msg_scheduler.mreg_6[26] ),
    .A2(_04474_),
    .B1(_04480_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00678_));
 sky130_fd_sc_hd__clkbuf_2 _10429_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04481_));
 sky130_fd_sc_hd__or2_1 _10430_ (.A(\sha256cu.msg_scheduler.mreg_7[27] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04482_));
 sky130_fd_sc_hd__o211a_1 _10431_ (.A1(\sha256cu.msg_scheduler.mreg_6[27] ),
    .A2(_04474_),
    .B1(_04482_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00679_));
 sky130_fd_sc_hd__or2_1 _10432_ (.A(\sha256cu.msg_scheduler.mreg_7[28] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04483_));
 sky130_fd_sc_hd__o211a_1 _10433_ (.A1(\sha256cu.msg_scheduler.mreg_6[28] ),
    .A2(_04474_),
    .B1(_04483_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00680_));
 sky130_fd_sc_hd__or2_1 _10434_ (.A(\sha256cu.msg_scheduler.mreg_7[29] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04484_));
 sky130_fd_sc_hd__o211a_1 _10435_ (.A1(\sha256cu.msg_scheduler.mreg_6[29] ),
    .A2(_04474_),
    .B1(_04484_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00681_));
 sky130_fd_sc_hd__or2_1 _10436_ (.A(\sha256cu.msg_scheduler.mreg_7[30] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04485_));
 sky130_fd_sc_hd__o211a_1 _10437_ (.A1(\sha256cu.msg_scheduler.mreg_6[30] ),
    .A2(_04474_),
    .B1(_04485_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00682_));
 sky130_fd_sc_hd__or2_1 _10438_ (.A(\sha256cu.msg_scheduler.mreg_7[31] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04486_));
 sky130_fd_sc_hd__o211a_1 _10439_ (.A1(\sha256cu.msg_scheduler.mreg_6[31] ),
    .A2(_04474_),
    .B1(_04486_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00683_));
 sky130_fd_sc_hd__buf_2 _10440_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04487_));
 sky130_fd_sc_hd__or2_1 _10441_ (.A(\sha256cu.msg_scheduler.mreg_8[0] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04488_));
 sky130_fd_sc_hd__o211a_1 _10442_ (.A1(\sha256cu.msg_scheduler.mreg_7[0] ),
    .A2(_04487_),
    .B1(_04488_),
    .C1(_04477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00684_));
 sky130_fd_sc_hd__or2_1 _10443_ (.A(\sha256cu.msg_scheduler.mreg_8[1] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04489_));
 sky130_fd_sc_hd__buf_2 _10444_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04490_));
 sky130_fd_sc_hd__o211a_1 _10445_ (.A1(\sha256cu.msg_scheduler.mreg_7[1] ),
    .A2(_04487_),
    .B1(_04489_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00685_));
 sky130_fd_sc_hd__or2_1 _10446_ (.A(\sha256cu.msg_scheduler.mreg_8[2] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04491_));
 sky130_fd_sc_hd__o211a_1 _10447_ (.A1(\sha256cu.msg_scheduler.mreg_7[2] ),
    .A2(_04487_),
    .B1(_04491_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00686_));
 sky130_fd_sc_hd__or2_1 _10448_ (.A(\sha256cu.msg_scheduler.mreg_8[3] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04492_));
 sky130_fd_sc_hd__o211a_1 _10449_ (.A1(\sha256cu.msg_scheduler.mreg_7[3] ),
    .A2(_04487_),
    .B1(_04492_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00687_));
 sky130_fd_sc_hd__or2_1 _10450_ (.A(\sha256cu.msg_scheduler.mreg_8[4] ),
    .B(_04481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04493_));
 sky130_fd_sc_hd__o211a_1 _10451_ (.A1(\sha256cu.msg_scheduler.mreg_7[4] ),
    .A2(_04487_),
    .B1(_04493_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00688_));
 sky130_fd_sc_hd__clkbuf_2 _10452_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04494_));
 sky130_fd_sc_hd__or2_1 _10453_ (.A(\sha256cu.msg_scheduler.mreg_8[5] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04495_));
 sky130_fd_sc_hd__o211a_1 _10454_ (.A1(\sha256cu.msg_scheduler.mreg_7[5] ),
    .A2(_04487_),
    .B1(_04495_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00689_));
 sky130_fd_sc_hd__or2_1 _10455_ (.A(\sha256cu.msg_scheduler.mreg_8[6] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04496_));
 sky130_fd_sc_hd__o211a_1 _10456_ (.A1(\sha256cu.msg_scheduler.mreg_7[6] ),
    .A2(_04487_),
    .B1(_04496_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00690_));
 sky130_fd_sc_hd__or2_1 _10457_ (.A(\sha256cu.msg_scheduler.mreg_8[7] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04497_));
 sky130_fd_sc_hd__o211a_1 _10458_ (.A1(\sha256cu.msg_scheduler.mreg_7[7] ),
    .A2(_04487_),
    .B1(_04497_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00691_));
 sky130_fd_sc_hd__or2_1 _10459_ (.A(\sha256cu.msg_scheduler.mreg_8[8] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04498_));
 sky130_fd_sc_hd__o211a_1 _10460_ (.A1(\sha256cu.msg_scheduler.mreg_7[8] ),
    .A2(_04487_),
    .B1(_04498_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00692_));
 sky130_fd_sc_hd__or2_1 _10461_ (.A(\sha256cu.msg_scheduler.mreg_8[9] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04499_));
 sky130_fd_sc_hd__o211a_1 _10462_ (.A1(\sha256cu.msg_scheduler.mreg_7[9] ),
    .A2(_04487_),
    .B1(_04499_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00693_));
 sky130_fd_sc_hd__clkbuf_4 _10463_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04500_));
 sky130_fd_sc_hd__or2_1 _10464_ (.A(\sha256cu.msg_scheduler.mreg_8[10] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04501_));
 sky130_fd_sc_hd__o211a_1 _10465_ (.A1(\sha256cu.msg_scheduler.mreg_7[10] ),
    .A2(_04500_),
    .B1(_04501_),
    .C1(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00694_));
 sky130_fd_sc_hd__or2_1 _10466_ (.A(\sha256cu.msg_scheduler.mreg_8[11] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04502_));
 sky130_fd_sc_hd__buf_2 _10467_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04503_));
 sky130_fd_sc_hd__o211a_1 _10468_ (.A1(\sha256cu.msg_scheduler.mreg_7[11] ),
    .A2(_04500_),
    .B1(_04502_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00695_));
 sky130_fd_sc_hd__or2_1 _10469_ (.A(\sha256cu.msg_scheduler.mreg_8[12] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04504_));
 sky130_fd_sc_hd__o211a_1 _10470_ (.A1(\sha256cu.msg_scheduler.mreg_7[12] ),
    .A2(_04500_),
    .B1(_04504_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00696_));
 sky130_fd_sc_hd__or2_1 _10471_ (.A(\sha256cu.msg_scheduler.mreg_8[13] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04505_));
 sky130_fd_sc_hd__o211a_1 _10472_ (.A1(\sha256cu.msg_scheduler.mreg_7[13] ),
    .A2(_04500_),
    .B1(_04505_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00697_));
 sky130_fd_sc_hd__or2_1 _10473_ (.A(\sha256cu.msg_scheduler.mreg_8[14] ),
    .B(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04506_));
 sky130_fd_sc_hd__o211a_1 _10474_ (.A1(\sha256cu.msg_scheduler.mreg_7[14] ),
    .A2(_04500_),
    .B1(_04506_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00698_));
 sky130_fd_sc_hd__clkbuf_2 _10475_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04507_));
 sky130_fd_sc_hd__or2_1 _10476_ (.A(\sha256cu.msg_scheduler.mreg_8[15] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04508_));
 sky130_fd_sc_hd__o211a_1 _10477_ (.A1(\sha256cu.msg_scheduler.mreg_7[15] ),
    .A2(_04500_),
    .B1(_04508_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00699_));
 sky130_fd_sc_hd__or2_1 _10478_ (.A(\sha256cu.msg_scheduler.mreg_8[16] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04509_));
 sky130_fd_sc_hd__o211a_1 _10479_ (.A1(\sha256cu.msg_scheduler.mreg_7[16] ),
    .A2(_04500_),
    .B1(_04509_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00700_));
 sky130_fd_sc_hd__or2_1 _10480_ (.A(\sha256cu.msg_scheduler.mreg_8[17] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04510_));
 sky130_fd_sc_hd__o211a_1 _10481_ (.A1(\sha256cu.msg_scheduler.mreg_7[17] ),
    .A2(_04500_),
    .B1(_04510_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00701_));
 sky130_fd_sc_hd__or2_1 _10482_ (.A(\sha256cu.msg_scheduler.mreg_8[18] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04511_));
 sky130_fd_sc_hd__o211a_1 _10483_ (.A1(\sha256cu.msg_scheduler.mreg_7[18] ),
    .A2(_04500_),
    .B1(_04511_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00702_));
 sky130_fd_sc_hd__or2_1 _10484_ (.A(\sha256cu.msg_scheduler.mreg_8[19] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04512_));
 sky130_fd_sc_hd__o211a_1 _10485_ (.A1(\sha256cu.msg_scheduler.mreg_7[19] ),
    .A2(_04500_),
    .B1(_04512_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00703_));
 sky130_fd_sc_hd__buf_2 _10486_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04513_));
 sky130_fd_sc_hd__or2_1 _10487_ (.A(\sha256cu.msg_scheduler.mreg_8[20] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04514_));
 sky130_fd_sc_hd__o211a_1 _10488_ (.A1(\sha256cu.msg_scheduler.mreg_7[20] ),
    .A2(_04513_),
    .B1(_04514_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00704_));
 sky130_fd_sc_hd__or2_1 _10489_ (.A(\sha256cu.msg_scheduler.mreg_8[21] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04515_));
 sky130_fd_sc_hd__buf_2 _10490_ (.A(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04516_));
 sky130_fd_sc_hd__o211a_1 _10491_ (.A1(\sha256cu.msg_scheduler.mreg_7[21] ),
    .A2(_04513_),
    .B1(_04515_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00705_));
 sky130_fd_sc_hd__or2_1 _10492_ (.A(\sha256cu.msg_scheduler.mreg_8[22] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04517_));
 sky130_fd_sc_hd__o211a_1 _10493_ (.A1(\sha256cu.msg_scheduler.mreg_7[22] ),
    .A2(_04513_),
    .B1(_04517_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00706_));
 sky130_fd_sc_hd__or2_1 _10494_ (.A(\sha256cu.msg_scheduler.mreg_8[23] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04518_));
 sky130_fd_sc_hd__o211a_1 _10495_ (.A1(\sha256cu.msg_scheduler.mreg_7[23] ),
    .A2(_04513_),
    .B1(_04518_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00707_));
 sky130_fd_sc_hd__or2_1 _10496_ (.A(\sha256cu.msg_scheduler.mreg_8[24] ),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04519_));
 sky130_fd_sc_hd__o211a_1 _10497_ (.A1(\sha256cu.msg_scheduler.mreg_7[24] ),
    .A2(_04513_),
    .B1(_04519_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00708_));
 sky130_fd_sc_hd__clkbuf_2 _10498_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04520_));
 sky130_fd_sc_hd__or2_1 _10499_ (.A(\sha256cu.msg_scheduler.mreg_8[25] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04521_));
 sky130_fd_sc_hd__o211a_1 _10500_ (.A1(\sha256cu.msg_scheduler.mreg_7[25] ),
    .A2(_04513_),
    .B1(_04521_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00709_));
 sky130_fd_sc_hd__or2_1 _10501_ (.A(\sha256cu.msg_scheduler.mreg_8[26] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04522_));
 sky130_fd_sc_hd__o211a_1 _10502_ (.A1(\sha256cu.msg_scheduler.mreg_7[26] ),
    .A2(_04513_),
    .B1(_04522_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00710_));
 sky130_fd_sc_hd__or2_1 _10503_ (.A(\sha256cu.msg_scheduler.mreg_8[27] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04523_));
 sky130_fd_sc_hd__o211a_1 _10504_ (.A1(\sha256cu.msg_scheduler.mreg_7[27] ),
    .A2(_04513_),
    .B1(_04523_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00711_));
 sky130_fd_sc_hd__or2_1 _10505_ (.A(\sha256cu.msg_scheduler.mreg_8[28] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04524_));
 sky130_fd_sc_hd__o211a_1 _10506_ (.A1(\sha256cu.msg_scheduler.mreg_7[28] ),
    .A2(_04513_),
    .B1(_04524_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00712_));
 sky130_fd_sc_hd__or2_1 _10507_ (.A(\sha256cu.msg_scheduler.mreg_8[29] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04525_));
 sky130_fd_sc_hd__o211a_1 _10508_ (.A1(\sha256cu.msg_scheduler.mreg_7[29] ),
    .A2(_04513_),
    .B1(_04525_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00713_));
 sky130_fd_sc_hd__buf_2 _10509_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04526_));
 sky130_fd_sc_hd__or2_1 _10510_ (.A(\sha256cu.msg_scheduler.mreg_8[30] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04527_));
 sky130_fd_sc_hd__o211a_1 _10511_ (.A1(\sha256cu.msg_scheduler.mreg_7[30] ),
    .A2(_04526_),
    .B1(_04527_),
    .C1(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00714_));
 sky130_fd_sc_hd__or2_1 _10512_ (.A(\sha256cu.msg_scheduler.mreg_8[31] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04528_));
 sky130_fd_sc_hd__buf_2 _10513_ (.A(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04529_));
 sky130_fd_sc_hd__buf_2 _10514_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04530_));
 sky130_fd_sc_hd__o211a_1 _10515_ (.A1(\sha256cu.msg_scheduler.mreg_7[31] ),
    .A2(_04526_),
    .B1(_04528_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00715_));
 sky130_fd_sc_hd__or2_1 _10516_ (.A(\sha256cu.msg_scheduler.mreg_9[0] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04531_));
 sky130_fd_sc_hd__o211a_1 _10517_ (.A1(\sha256cu.msg_scheduler.mreg_8[0] ),
    .A2(_04526_),
    .B1(_04531_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00716_));
 sky130_fd_sc_hd__or2_1 _10518_ (.A(\sha256cu.msg_scheduler.mreg_9[1] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04532_));
 sky130_fd_sc_hd__o211a_1 _10519_ (.A1(\sha256cu.msg_scheduler.mreg_8[1] ),
    .A2(_04526_),
    .B1(_04532_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00717_));
 sky130_fd_sc_hd__or2_1 _10520_ (.A(\sha256cu.msg_scheduler.mreg_9[2] ),
    .B(_04520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04533_));
 sky130_fd_sc_hd__o211a_1 _10521_ (.A1(\sha256cu.msg_scheduler.mreg_8[2] ),
    .A2(_04526_),
    .B1(_04533_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00718_));
 sky130_fd_sc_hd__clkbuf_2 _10522_ (.A(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04534_));
 sky130_fd_sc_hd__or2_1 _10523_ (.A(\sha256cu.msg_scheduler.mreg_9[3] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04535_));
 sky130_fd_sc_hd__o211a_1 _10524_ (.A1(\sha256cu.msg_scheduler.mreg_8[3] ),
    .A2(_04526_),
    .B1(_04535_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00719_));
 sky130_fd_sc_hd__or2_1 _10525_ (.A(\sha256cu.msg_scheduler.mreg_9[4] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04536_));
 sky130_fd_sc_hd__o211a_1 _10526_ (.A1(\sha256cu.msg_scheduler.mreg_8[4] ),
    .A2(_04526_),
    .B1(_04536_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00720_));
 sky130_fd_sc_hd__or2_1 _10527_ (.A(\sha256cu.msg_scheduler.mreg_9[5] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04537_));
 sky130_fd_sc_hd__o211a_1 _10528_ (.A1(\sha256cu.msg_scheduler.mreg_8[5] ),
    .A2(_04526_),
    .B1(_04537_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00721_));
 sky130_fd_sc_hd__or2_1 _10529_ (.A(\sha256cu.msg_scheduler.mreg_9[6] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04538_));
 sky130_fd_sc_hd__o211a_1 _10530_ (.A1(\sha256cu.msg_scheduler.mreg_8[6] ),
    .A2(_04526_),
    .B1(_04538_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00722_));
 sky130_fd_sc_hd__or2_1 _10531_ (.A(\sha256cu.msg_scheduler.mreg_9[7] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04539_));
 sky130_fd_sc_hd__o211a_1 _10532_ (.A1(\sha256cu.msg_scheduler.mreg_8[7] ),
    .A2(_04526_),
    .B1(_04539_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00723_));
 sky130_fd_sc_hd__buf_2 _10533_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04540_));
 sky130_fd_sc_hd__or2_1 _10534_ (.A(\sha256cu.msg_scheduler.mreg_9[8] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04541_));
 sky130_fd_sc_hd__o211a_1 _10535_ (.A1(\sha256cu.msg_scheduler.mreg_8[8] ),
    .A2(_04540_),
    .B1(_04541_),
    .C1(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00724_));
 sky130_fd_sc_hd__or2_1 _10536_ (.A(\sha256cu.msg_scheduler.mreg_9[9] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04542_));
 sky130_fd_sc_hd__buf_2 _10537_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04543_));
 sky130_fd_sc_hd__o211a_1 _10538_ (.A1(\sha256cu.msg_scheduler.mreg_8[9] ),
    .A2(_04540_),
    .B1(_04542_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00725_));
 sky130_fd_sc_hd__or2_1 _10539_ (.A(\sha256cu.msg_scheduler.mreg_9[10] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04544_));
 sky130_fd_sc_hd__o211a_1 _10540_ (.A1(\sha256cu.msg_scheduler.mreg_8[10] ),
    .A2(_04540_),
    .B1(_04544_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00726_));
 sky130_fd_sc_hd__or2_1 _10541_ (.A(\sha256cu.msg_scheduler.mreg_9[11] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04545_));
 sky130_fd_sc_hd__o211a_1 _10542_ (.A1(\sha256cu.msg_scheduler.mreg_8[11] ),
    .A2(_04540_),
    .B1(_04545_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00727_));
 sky130_fd_sc_hd__or2_1 _10543_ (.A(\sha256cu.msg_scheduler.mreg_9[12] ),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04546_));
 sky130_fd_sc_hd__o211a_1 _10544_ (.A1(\sha256cu.msg_scheduler.mreg_8[12] ),
    .A2(_04540_),
    .B1(_04546_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00728_));
 sky130_fd_sc_hd__clkbuf_4 _10545_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04547_));
 sky130_fd_sc_hd__clkbuf_2 _10546_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04548_));
 sky130_fd_sc_hd__or2_1 _10547_ (.A(\sha256cu.msg_scheduler.mreg_9[13] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04549_));
 sky130_fd_sc_hd__o211a_1 _10548_ (.A1(\sha256cu.msg_scheduler.mreg_8[13] ),
    .A2(_04540_),
    .B1(_04549_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00729_));
 sky130_fd_sc_hd__or2_1 _10549_ (.A(\sha256cu.msg_scheduler.mreg_9[14] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04550_));
 sky130_fd_sc_hd__o211a_1 _10550_ (.A1(\sha256cu.msg_scheduler.mreg_8[14] ),
    .A2(_04540_),
    .B1(_04550_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00730_));
 sky130_fd_sc_hd__or2_1 _10551_ (.A(\sha256cu.msg_scheduler.mreg_9[15] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04551_));
 sky130_fd_sc_hd__o211a_1 _10552_ (.A1(\sha256cu.msg_scheduler.mreg_8[15] ),
    .A2(_04540_),
    .B1(_04551_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00731_));
 sky130_fd_sc_hd__or2_1 _10553_ (.A(\sha256cu.msg_scheduler.mreg_9[16] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04552_));
 sky130_fd_sc_hd__o211a_1 _10554_ (.A1(\sha256cu.msg_scheduler.mreg_8[16] ),
    .A2(_04540_),
    .B1(_04552_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00732_));
 sky130_fd_sc_hd__or2_1 _10555_ (.A(\sha256cu.msg_scheduler.mreg_9[17] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04553_));
 sky130_fd_sc_hd__o211a_1 _10556_ (.A1(\sha256cu.msg_scheduler.mreg_8[17] ),
    .A2(_04540_),
    .B1(_04553_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00733_));
 sky130_fd_sc_hd__buf_2 _10557_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04554_));
 sky130_fd_sc_hd__or2_1 _10558_ (.A(\sha256cu.msg_scheduler.mreg_9[18] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04555_));
 sky130_fd_sc_hd__o211a_1 _10559_ (.A1(\sha256cu.msg_scheduler.mreg_8[18] ),
    .A2(_04554_),
    .B1(_04555_),
    .C1(_04543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _10560_ (.A(\sha256cu.msg_scheduler.mreg_9[19] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04556_));
 sky130_fd_sc_hd__buf_2 _10561_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04557_));
 sky130_fd_sc_hd__o211a_1 _10562_ (.A1(\sha256cu.msg_scheduler.mreg_8[19] ),
    .A2(_04554_),
    .B1(_04556_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00735_));
 sky130_fd_sc_hd__or2_1 _10563_ (.A(\sha256cu.msg_scheduler.mreg_9[20] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04558_));
 sky130_fd_sc_hd__o211a_1 _10564_ (.A1(\sha256cu.msg_scheduler.mreg_8[20] ),
    .A2(_04554_),
    .B1(_04558_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _10565_ (.A(\sha256cu.msg_scheduler.mreg_9[21] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04559_));
 sky130_fd_sc_hd__o211a_1 _10566_ (.A1(\sha256cu.msg_scheduler.mreg_8[21] ),
    .A2(_04554_),
    .B1(_04559_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00737_));
 sky130_fd_sc_hd__or2_1 _10567_ (.A(\sha256cu.msg_scheduler.mreg_9[22] ),
    .B(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04560_));
 sky130_fd_sc_hd__o211a_1 _10568_ (.A1(\sha256cu.msg_scheduler.mreg_8[22] ),
    .A2(_04554_),
    .B1(_04560_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00738_));
 sky130_fd_sc_hd__clkbuf_2 _10569_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04561_));
 sky130_fd_sc_hd__or2_1 _10570_ (.A(\sha256cu.msg_scheduler.mreg_9[23] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04562_));
 sky130_fd_sc_hd__o211a_1 _10571_ (.A1(\sha256cu.msg_scheduler.mreg_8[23] ),
    .A2(_04554_),
    .B1(_04562_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00739_));
 sky130_fd_sc_hd__or2_1 _10572_ (.A(\sha256cu.msg_scheduler.mreg_9[24] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04563_));
 sky130_fd_sc_hd__o211a_1 _10573_ (.A1(\sha256cu.msg_scheduler.mreg_8[24] ),
    .A2(_04554_),
    .B1(_04563_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00740_));
 sky130_fd_sc_hd__or2_1 _10574_ (.A(\sha256cu.msg_scheduler.mreg_9[25] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04564_));
 sky130_fd_sc_hd__o211a_1 _10575_ (.A1(\sha256cu.msg_scheduler.mreg_8[25] ),
    .A2(_04554_),
    .B1(_04564_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00741_));
 sky130_fd_sc_hd__or2_1 _10576_ (.A(\sha256cu.msg_scheduler.mreg_9[26] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04565_));
 sky130_fd_sc_hd__o211a_1 _10577_ (.A1(\sha256cu.msg_scheduler.mreg_8[26] ),
    .A2(_04554_),
    .B1(_04565_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00742_));
 sky130_fd_sc_hd__or2_1 _10578_ (.A(\sha256cu.msg_scheduler.mreg_9[27] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04566_));
 sky130_fd_sc_hd__o211a_1 _10579_ (.A1(\sha256cu.msg_scheduler.mreg_8[27] ),
    .A2(_04554_),
    .B1(_04566_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00743_));
 sky130_fd_sc_hd__buf_2 _10580_ (.A(_04447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04567_));
 sky130_fd_sc_hd__or2_1 _10581_ (.A(\sha256cu.msg_scheduler.mreg_9[28] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04568_));
 sky130_fd_sc_hd__o211a_1 _10582_ (.A1(\sha256cu.msg_scheduler.mreg_8[28] ),
    .A2(_04567_),
    .B1(_04568_),
    .C1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00744_));
 sky130_fd_sc_hd__or2_1 _10583_ (.A(\sha256cu.msg_scheduler.mreg_9[29] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04569_));
 sky130_fd_sc_hd__buf_2 _10584_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04570_));
 sky130_fd_sc_hd__o211a_1 _10585_ (.A1(\sha256cu.msg_scheduler.mreg_8[29] ),
    .A2(_04567_),
    .B1(_04569_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _10586_ (.A(\sha256cu.msg_scheduler.mreg_9[30] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04571_));
 sky130_fd_sc_hd__o211a_1 _10587_ (.A1(\sha256cu.msg_scheduler.mreg_8[30] ),
    .A2(_04567_),
    .B1(_04571_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00746_));
 sky130_fd_sc_hd__or2_1 _10588_ (.A(\sha256cu.msg_scheduler.mreg_9[31] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04572_));
 sky130_fd_sc_hd__o211a_1 _10589_ (.A1(\sha256cu.msg_scheduler.mreg_8[31] ),
    .A2(_04567_),
    .B1(_04572_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00747_));
 sky130_fd_sc_hd__or2_1 _10590_ (.A(\sha256cu.msg_scheduler.mreg_10[0] ),
    .B(_04561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04573_));
 sky130_fd_sc_hd__o211a_1 _10591_ (.A1(\sha256cu.msg_scheduler.mreg_9[0] ),
    .A2(_04567_),
    .B1(_04573_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00748_));
 sky130_fd_sc_hd__clkbuf_2 _10592_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04574_));
 sky130_fd_sc_hd__or2_1 _10593_ (.A(\sha256cu.msg_scheduler.mreg_10[1] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04575_));
 sky130_fd_sc_hd__o211a_1 _10594_ (.A1(\sha256cu.msg_scheduler.mreg_9[1] ),
    .A2(_04567_),
    .B1(_04575_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00749_));
 sky130_fd_sc_hd__or2_1 _10595_ (.A(\sha256cu.msg_scheduler.mreg_10[2] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04576_));
 sky130_fd_sc_hd__o211a_1 _10596_ (.A1(\sha256cu.msg_scheduler.mreg_9[2] ),
    .A2(_04567_),
    .B1(_04576_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00750_));
 sky130_fd_sc_hd__or2_1 _10597_ (.A(\sha256cu.msg_scheduler.mreg_10[3] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04577_));
 sky130_fd_sc_hd__o211a_1 _10598_ (.A1(\sha256cu.msg_scheduler.mreg_9[3] ),
    .A2(_04567_),
    .B1(_04577_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00751_));
 sky130_fd_sc_hd__or2_1 _10599_ (.A(\sha256cu.msg_scheduler.mreg_10[4] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04578_));
 sky130_fd_sc_hd__o211a_1 _10600_ (.A1(\sha256cu.msg_scheduler.mreg_9[4] ),
    .A2(_04567_),
    .B1(_04578_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00752_));
 sky130_fd_sc_hd__or2_1 _10601_ (.A(\sha256cu.msg_scheduler.mreg_10[5] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04579_));
 sky130_fd_sc_hd__o211a_1 _10602_ (.A1(\sha256cu.msg_scheduler.mreg_9[5] ),
    .A2(_04567_),
    .B1(_04579_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00753_));
 sky130_fd_sc_hd__clkbuf_4 _10603_ (.A(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04580_));
 sky130_fd_sc_hd__clkbuf_4 _10604_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04581_));
 sky130_fd_sc_hd__or2_1 _10605_ (.A(\sha256cu.msg_scheduler.mreg_10[6] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04582_));
 sky130_fd_sc_hd__o211a_1 _10606_ (.A1(\sha256cu.msg_scheduler.mreg_9[6] ),
    .A2(_04581_),
    .B1(_04582_),
    .C1(_04570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00754_));
 sky130_fd_sc_hd__or2_1 _10607_ (.A(\sha256cu.msg_scheduler.mreg_10[7] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04583_));
 sky130_fd_sc_hd__buf_2 _10608_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04584_));
 sky130_fd_sc_hd__o211a_1 _10609_ (.A1(\sha256cu.msg_scheduler.mreg_9[7] ),
    .A2(_04581_),
    .B1(_04583_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00755_));
 sky130_fd_sc_hd__or2_1 _10610_ (.A(\sha256cu.msg_scheduler.mreg_10[8] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04585_));
 sky130_fd_sc_hd__o211a_1 _10611_ (.A1(\sha256cu.msg_scheduler.mreg_9[8] ),
    .A2(_04581_),
    .B1(_04585_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _10612_ (.A(\sha256cu.msg_scheduler.mreg_10[9] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04586_));
 sky130_fd_sc_hd__o211a_1 _10613_ (.A1(\sha256cu.msg_scheduler.mreg_9[9] ),
    .A2(_04581_),
    .B1(_04586_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _10614_ (.A(\sha256cu.msg_scheduler.mreg_10[10] ),
    .B(_04574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04587_));
 sky130_fd_sc_hd__o211a_1 _10615_ (.A1(\sha256cu.msg_scheduler.mreg_9[10] ),
    .A2(_04581_),
    .B1(_04587_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00758_));
 sky130_fd_sc_hd__clkbuf_2 _10616_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04588_));
 sky130_fd_sc_hd__or2_1 _10617_ (.A(\sha256cu.msg_scheduler.mreg_10[11] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04589_));
 sky130_fd_sc_hd__o211a_1 _10618_ (.A1(\sha256cu.msg_scheduler.mreg_9[11] ),
    .A2(_04581_),
    .B1(_04589_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _10619_ (.A(\sha256cu.msg_scheduler.mreg_10[12] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04590_));
 sky130_fd_sc_hd__o211a_1 _10620_ (.A1(\sha256cu.msg_scheduler.mreg_9[12] ),
    .A2(_04581_),
    .B1(_04590_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _10621_ (.A(\sha256cu.msg_scheduler.mreg_10[13] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04591_));
 sky130_fd_sc_hd__o211a_1 _10622_ (.A1(\sha256cu.msg_scheduler.mreg_9[13] ),
    .A2(_04581_),
    .B1(_04591_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _10623_ (.A(\sha256cu.msg_scheduler.mreg_10[14] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04592_));
 sky130_fd_sc_hd__o211a_1 _10624_ (.A1(\sha256cu.msg_scheduler.mreg_9[14] ),
    .A2(_04581_),
    .B1(_04592_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _10625_ (.A(\sha256cu.msg_scheduler.mreg_10[15] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04593_));
 sky130_fd_sc_hd__o211a_1 _10626_ (.A1(\sha256cu.msg_scheduler.mreg_9[15] ),
    .A2(_04581_),
    .B1(_04593_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00763_));
 sky130_fd_sc_hd__buf_2 _10627_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04594_));
 sky130_fd_sc_hd__or2_1 _10628_ (.A(\sha256cu.msg_scheduler.mreg_10[16] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04595_));
 sky130_fd_sc_hd__o211a_1 _10629_ (.A1(\sha256cu.msg_scheduler.mreg_9[16] ),
    .A2(_04594_),
    .B1(_04595_),
    .C1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _10630_ (.A(\sha256cu.msg_scheduler.mreg_10[17] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04596_));
 sky130_fd_sc_hd__buf_2 _10631_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04597_));
 sky130_fd_sc_hd__o211a_1 _10632_ (.A1(\sha256cu.msg_scheduler.mreg_9[17] ),
    .A2(_04594_),
    .B1(_04596_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _10633_ (.A(\sha256cu.msg_scheduler.mreg_10[18] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04598_));
 sky130_fd_sc_hd__o211a_1 _10634_ (.A1(\sha256cu.msg_scheduler.mreg_9[18] ),
    .A2(_04594_),
    .B1(_04598_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00766_));
 sky130_fd_sc_hd__or2_1 _10635_ (.A(\sha256cu.msg_scheduler.mreg_10[19] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04599_));
 sky130_fd_sc_hd__o211a_1 _10636_ (.A1(\sha256cu.msg_scheduler.mreg_9[19] ),
    .A2(_04594_),
    .B1(_04599_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _10637_ (.A(\sha256cu.msg_scheduler.mreg_10[20] ),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04600_));
 sky130_fd_sc_hd__o211a_1 _10638_ (.A1(\sha256cu.msg_scheduler.mreg_9[20] ),
    .A2(_04594_),
    .B1(_04600_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00768_));
 sky130_fd_sc_hd__clkbuf_2 _10639_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04601_));
 sky130_fd_sc_hd__or2_1 _10640_ (.A(\sha256cu.msg_scheduler.mreg_10[21] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04602_));
 sky130_fd_sc_hd__o211a_1 _10641_ (.A1(\sha256cu.msg_scheduler.mreg_9[21] ),
    .A2(_04594_),
    .B1(_04602_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _10642_ (.A(\sha256cu.msg_scheduler.mreg_10[22] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04603_));
 sky130_fd_sc_hd__o211a_1 _10643_ (.A1(\sha256cu.msg_scheduler.mreg_9[22] ),
    .A2(_04594_),
    .B1(_04603_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00770_));
 sky130_fd_sc_hd__or2_1 _10644_ (.A(\sha256cu.msg_scheduler.mreg_10[23] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04604_));
 sky130_fd_sc_hd__o211a_1 _10645_ (.A1(\sha256cu.msg_scheduler.mreg_9[23] ),
    .A2(_04594_),
    .B1(_04604_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _10646_ (.A(\sha256cu.msg_scheduler.mreg_10[24] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04605_));
 sky130_fd_sc_hd__o211a_1 _10647_ (.A1(\sha256cu.msg_scheduler.mreg_9[24] ),
    .A2(_04594_),
    .B1(_04605_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _10648_ (.A(\sha256cu.msg_scheduler.mreg_10[25] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04606_));
 sky130_fd_sc_hd__o211a_1 _10649_ (.A1(\sha256cu.msg_scheduler.mreg_9[25] ),
    .A2(_04594_),
    .B1(_04606_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00773_));
 sky130_fd_sc_hd__buf_2 _10650_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04607_));
 sky130_fd_sc_hd__or2_1 _10651_ (.A(\sha256cu.msg_scheduler.mreg_10[26] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04608_));
 sky130_fd_sc_hd__o211a_1 _10652_ (.A1(\sha256cu.msg_scheduler.mreg_9[26] ),
    .A2(_04607_),
    .B1(_04608_),
    .C1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _10653_ (.A(\sha256cu.msg_scheduler.mreg_10[27] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04609_));
 sky130_fd_sc_hd__buf_2 _10654_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04610_));
 sky130_fd_sc_hd__o211a_1 _10655_ (.A1(\sha256cu.msg_scheduler.mreg_9[27] ),
    .A2(_04607_),
    .B1(_04609_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _10656_ (.A(\sha256cu.msg_scheduler.mreg_10[28] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04611_));
 sky130_fd_sc_hd__o211a_1 _10657_ (.A1(\sha256cu.msg_scheduler.mreg_9[28] ),
    .A2(_04607_),
    .B1(_04611_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _10658_ (.A(\sha256cu.msg_scheduler.mreg_10[29] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04612_));
 sky130_fd_sc_hd__o211a_1 _10659_ (.A1(\sha256cu.msg_scheduler.mreg_9[29] ),
    .A2(_04607_),
    .B1(_04612_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _10660_ (.A(\sha256cu.msg_scheduler.mreg_10[30] ),
    .B(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04613_));
 sky130_fd_sc_hd__o211a_1 _10661_ (.A1(\sha256cu.msg_scheduler.mreg_9[30] ),
    .A2(_04607_),
    .B1(_04613_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00778_));
 sky130_fd_sc_hd__clkbuf_2 _10662_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04614_));
 sky130_fd_sc_hd__or2_1 _10663_ (.A(\sha256cu.msg_scheduler.mreg_10[31] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04615_));
 sky130_fd_sc_hd__o211a_1 _10664_ (.A1(\sha256cu.msg_scheduler.mreg_9[31] ),
    .A2(_04607_),
    .B1(_04615_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00779_));
 sky130_fd_sc_hd__or2_1 _10665_ (.A(\sha256cu.msg_scheduler.mreg_11[0] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04616_));
 sky130_fd_sc_hd__o211a_1 _10666_ (.A1(\sha256cu.msg_scheduler.mreg_10[0] ),
    .A2(_04607_),
    .B1(_04616_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00780_));
 sky130_fd_sc_hd__or2_1 _10667_ (.A(\sha256cu.msg_scheduler.mreg_11[1] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04617_));
 sky130_fd_sc_hd__o211a_1 _10668_ (.A1(\sha256cu.msg_scheduler.mreg_10[1] ),
    .A2(_04607_),
    .B1(_04617_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _10669_ (.A(\sha256cu.msg_scheduler.mreg_11[2] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04618_));
 sky130_fd_sc_hd__o211a_1 _10670_ (.A1(\sha256cu.msg_scheduler.mreg_10[2] ),
    .A2(_04607_),
    .B1(_04618_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00782_));
 sky130_fd_sc_hd__or2_1 _10671_ (.A(\sha256cu.msg_scheduler.mreg_11[3] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04619_));
 sky130_fd_sc_hd__o211a_1 _10672_ (.A1(\sha256cu.msg_scheduler.mreg_10[3] ),
    .A2(_04607_),
    .B1(_04619_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00783_));
 sky130_fd_sc_hd__buf_2 _10673_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04620_));
 sky130_fd_sc_hd__or2_1 _10674_ (.A(\sha256cu.msg_scheduler.mreg_11[4] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04621_));
 sky130_fd_sc_hd__o211a_1 _10675_ (.A1(\sha256cu.msg_scheduler.mreg_10[4] ),
    .A2(_04620_),
    .B1(_04621_),
    .C1(_04610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _10676_ (.A(\sha256cu.msg_scheduler.mreg_11[5] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04622_));
 sky130_fd_sc_hd__clkbuf_4 _10677_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04623_));
 sky130_fd_sc_hd__o211a_1 _10678_ (.A1(\sha256cu.msg_scheduler.mreg_10[5] ),
    .A2(_04620_),
    .B1(_04622_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00785_));
 sky130_fd_sc_hd__or2_1 _10679_ (.A(\sha256cu.msg_scheduler.mreg_11[6] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04624_));
 sky130_fd_sc_hd__o211a_1 _10680_ (.A1(\sha256cu.msg_scheduler.mreg_10[6] ),
    .A2(_04620_),
    .B1(_04624_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00786_));
 sky130_fd_sc_hd__or2_1 _10681_ (.A(\sha256cu.msg_scheduler.mreg_11[7] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04625_));
 sky130_fd_sc_hd__o211a_1 _10682_ (.A1(\sha256cu.msg_scheduler.mreg_10[7] ),
    .A2(_04620_),
    .B1(_04625_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00787_));
 sky130_fd_sc_hd__or2_1 _10683_ (.A(\sha256cu.msg_scheduler.mreg_11[8] ),
    .B(_04614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04626_));
 sky130_fd_sc_hd__o211a_1 _10684_ (.A1(\sha256cu.msg_scheduler.mreg_10[8] ),
    .A2(_04620_),
    .B1(_04626_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00788_));
 sky130_fd_sc_hd__clkbuf_2 _10685_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04627_));
 sky130_fd_sc_hd__or2_1 _10686_ (.A(\sha256cu.msg_scheduler.mreg_11[9] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04628_));
 sky130_fd_sc_hd__o211a_1 _10687_ (.A1(\sha256cu.msg_scheduler.mreg_10[9] ),
    .A2(_04620_),
    .B1(_04628_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00789_));
 sky130_fd_sc_hd__or2_1 _10688_ (.A(\sha256cu.msg_scheduler.mreg_11[10] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04629_));
 sky130_fd_sc_hd__o211a_1 _10689_ (.A1(\sha256cu.msg_scheduler.mreg_10[10] ),
    .A2(_04620_),
    .B1(_04629_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00790_));
 sky130_fd_sc_hd__or2_1 _10690_ (.A(\sha256cu.msg_scheduler.mreg_11[11] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04630_));
 sky130_fd_sc_hd__o211a_1 _10691_ (.A1(\sha256cu.msg_scheduler.mreg_10[11] ),
    .A2(_04620_),
    .B1(_04630_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00791_));
 sky130_fd_sc_hd__or2_1 _10692_ (.A(\sha256cu.msg_scheduler.mreg_11[12] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04631_));
 sky130_fd_sc_hd__o211a_1 _10693_ (.A1(\sha256cu.msg_scheduler.mreg_10[12] ),
    .A2(_04620_),
    .B1(_04631_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00792_));
 sky130_fd_sc_hd__or2_1 _10694_ (.A(\sha256cu.msg_scheduler.mreg_11[13] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04632_));
 sky130_fd_sc_hd__o211a_1 _10695_ (.A1(\sha256cu.msg_scheduler.mreg_10[13] ),
    .A2(_04620_),
    .B1(_04632_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00793_));
 sky130_fd_sc_hd__buf_2 _10696_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04633_));
 sky130_fd_sc_hd__or2_1 _10697_ (.A(\sha256cu.msg_scheduler.mreg_11[14] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04634_));
 sky130_fd_sc_hd__o211a_1 _10698_ (.A1(\sha256cu.msg_scheduler.mreg_10[14] ),
    .A2(_04633_),
    .B1(_04634_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _10699_ (.A(\sha256cu.msg_scheduler.mreg_11[15] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04635_));
 sky130_fd_sc_hd__buf_2 _10700_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04636_));
 sky130_fd_sc_hd__o211a_1 _10701_ (.A1(\sha256cu.msg_scheduler.mreg_10[15] ),
    .A2(_04633_),
    .B1(_04635_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _10702_ (.A(\sha256cu.msg_scheduler.mreg_11[16] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04637_));
 sky130_fd_sc_hd__o211a_1 _10703_ (.A1(\sha256cu.msg_scheduler.mreg_10[16] ),
    .A2(_04633_),
    .B1(_04637_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _10704_ (.A(\sha256cu.msg_scheduler.mreg_11[17] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04638_));
 sky130_fd_sc_hd__o211a_1 _10705_ (.A1(\sha256cu.msg_scheduler.mreg_10[17] ),
    .A2(_04633_),
    .B1(_04638_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _10706_ (.A(\sha256cu.msg_scheduler.mreg_11[18] ),
    .B(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04639_));
 sky130_fd_sc_hd__o211a_1 _10707_ (.A1(\sha256cu.msg_scheduler.mreg_10[18] ),
    .A2(_04633_),
    .B1(_04639_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00798_));
 sky130_fd_sc_hd__clkbuf_2 _10708_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04640_));
 sky130_fd_sc_hd__or2_1 _10709_ (.A(\sha256cu.msg_scheduler.mreg_11[19] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04641_));
 sky130_fd_sc_hd__o211a_1 _10710_ (.A1(\sha256cu.msg_scheduler.mreg_10[19] ),
    .A2(_04633_),
    .B1(_04641_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _10711_ (.A(\sha256cu.msg_scheduler.mreg_11[20] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04642_));
 sky130_fd_sc_hd__o211a_1 _10712_ (.A1(\sha256cu.msg_scheduler.mreg_10[20] ),
    .A2(_04633_),
    .B1(_04642_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00800_));
 sky130_fd_sc_hd__or2_1 _10713_ (.A(\sha256cu.msg_scheduler.mreg_11[21] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04643_));
 sky130_fd_sc_hd__o211a_1 _10714_ (.A1(\sha256cu.msg_scheduler.mreg_10[21] ),
    .A2(_04633_),
    .B1(_04643_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00801_));
 sky130_fd_sc_hd__or2_1 _10715_ (.A(\sha256cu.msg_scheduler.mreg_11[22] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04644_));
 sky130_fd_sc_hd__o211a_1 _10716_ (.A1(\sha256cu.msg_scheduler.mreg_10[22] ),
    .A2(_04633_),
    .B1(_04644_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _10717_ (.A(\sha256cu.msg_scheduler.mreg_11[23] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04645_));
 sky130_fd_sc_hd__o211a_1 _10718_ (.A1(\sha256cu.msg_scheduler.mreg_10[23] ),
    .A2(_04633_),
    .B1(_04645_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00803_));
 sky130_fd_sc_hd__clkbuf_4 _10719_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04646_));
 sky130_fd_sc_hd__or2_1 _10720_ (.A(\sha256cu.msg_scheduler.mreg_11[24] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04647_));
 sky130_fd_sc_hd__o211a_1 _10721_ (.A1(\sha256cu.msg_scheduler.mreg_10[24] ),
    .A2(_04646_),
    .B1(_04647_),
    .C1(_04636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00804_));
 sky130_fd_sc_hd__or2_1 _10722_ (.A(\sha256cu.msg_scheduler.mreg_11[25] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04648_));
 sky130_fd_sc_hd__buf_2 _10723_ (.A(_04529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04649_));
 sky130_fd_sc_hd__o211a_1 _10724_ (.A1(\sha256cu.msg_scheduler.mreg_10[25] ),
    .A2(_04646_),
    .B1(_04648_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _10725_ (.A(\sha256cu.msg_scheduler.mreg_11[26] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04650_));
 sky130_fd_sc_hd__o211a_1 _10726_ (.A1(\sha256cu.msg_scheduler.mreg_10[26] ),
    .A2(_04646_),
    .B1(_04650_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00806_));
 sky130_fd_sc_hd__or2_1 _10727_ (.A(\sha256cu.msg_scheduler.mreg_11[27] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04651_));
 sky130_fd_sc_hd__o211a_1 _10728_ (.A1(\sha256cu.msg_scheduler.mreg_10[27] ),
    .A2(_04646_),
    .B1(_04651_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _10729_ (.A(\sha256cu.msg_scheduler.mreg_11[28] ),
    .B(_04640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04652_));
 sky130_fd_sc_hd__o211a_1 _10730_ (.A1(\sha256cu.msg_scheduler.mreg_10[28] ),
    .A2(_04646_),
    .B1(_04652_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00808_));
 sky130_fd_sc_hd__clkbuf_2 _10731_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04653_));
 sky130_fd_sc_hd__or2_1 _10732_ (.A(\sha256cu.msg_scheduler.mreg_11[29] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04654_));
 sky130_fd_sc_hd__o211a_1 _10733_ (.A1(\sha256cu.msg_scheduler.mreg_10[29] ),
    .A2(_04646_),
    .B1(_04654_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _10734_ (.A(\sha256cu.msg_scheduler.mreg_11[30] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04655_));
 sky130_fd_sc_hd__o211a_1 _10735_ (.A1(\sha256cu.msg_scheduler.mreg_10[30] ),
    .A2(_04646_),
    .B1(_04655_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00810_));
 sky130_fd_sc_hd__or2_1 _10736_ (.A(\sha256cu.msg_scheduler.mreg_11[31] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04656_));
 sky130_fd_sc_hd__o211a_1 _10737_ (.A1(\sha256cu.msg_scheduler.mreg_10[31] ),
    .A2(_04646_),
    .B1(_04656_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _10738_ (.A(\sha256cu.msg_scheduler.mreg_12[0] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04657_));
 sky130_fd_sc_hd__o211a_1 _10739_ (.A1(\sha256cu.msg_scheduler.mreg_11[0] ),
    .A2(_04646_),
    .B1(_04657_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _10740_ (.A(\sha256cu.msg_scheduler.mreg_12[1] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04658_));
 sky130_fd_sc_hd__o211a_1 _10741_ (.A1(\sha256cu.msg_scheduler.mreg_11[1] ),
    .A2(_04646_),
    .B1(_04658_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00813_));
 sky130_fd_sc_hd__clkbuf_4 _10742_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04659_));
 sky130_fd_sc_hd__or2_1 _10743_ (.A(\sha256cu.msg_scheduler.mreg_12[2] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04660_));
 sky130_fd_sc_hd__o211a_1 _10744_ (.A1(\sha256cu.msg_scheduler.mreg_11[2] ),
    .A2(_04659_),
    .B1(_04660_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00814_));
 sky130_fd_sc_hd__or2_1 _10745_ (.A(\sha256cu.msg_scheduler.mreg_12[3] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_4 _10746_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04662_));
 sky130_fd_sc_hd__o211a_1 _10747_ (.A1(\sha256cu.msg_scheduler.mreg_11[3] ),
    .A2(_04659_),
    .B1(_04661_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00815_));
 sky130_fd_sc_hd__or2_1 _10748_ (.A(\sha256cu.msg_scheduler.mreg_12[4] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04663_));
 sky130_fd_sc_hd__o211a_1 _10749_ (.A1(\sha256cu.msg_scheduler.mreg_11[4] ),
    .A2(_04659_),
    .B1(_04663_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00816_));
 sky130_fd_sc_hd__or2_1 _10750_ (.A(\sha256cu.msg_scheduler.mreg_12[5] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04664_));
 sky130_fd_sc_hd__o211a_1 _10751_ (.A1(\sha256cu.msg_scheduler.mreg_11[5] ),
    .A2(_04659_),
    .B1(_04664_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _10752_ (.A(\sha256cu.msg_scheduler.mreg_12[6] ),
    .B(_04653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04665_));
 sky130_fd_sc_hd__o211a_1 _10753_ (.A1(\sha256cu.msg_scheduler.mreg_11[6] ),
    .A2(_04659_),
    .B1(_04665_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00818_));
 sky130_fd_sc_hd__clkbuf_2 _10754_ (.A(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04666_));
 sky130_fd_sc_hd__or2_1 _10755_ (.A(\sha256cu.msg_scheduler.mreg_12[7] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04667_));
 sky130_fd_sc_hd__o211a_1 _10756_ (.A1(\sha256cu.msg_scheduler.mreg_11[7] ),
    .A2(_04659_),
    .B1(_04667_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00819_));
 sky130_fd_sc_hd__or2_1 _10757_ (.A(\sha256cu.msg_scheduler.mreg_12[8] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04668_));
 sky130_fd_sc_hd__o211a_1 _10758_ (.A1(\sha256cu.msg_scheduler.mreg_11[8] ),
    .A2(_04659_),
    .B1(_04668_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00820_));
 sky130_fd_sc_hd__or2_1 _10759_ (.A(\sha256cu.msg_scheduler.mreg_12[9] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04669_));
 sky130_fd_sc_hd__o211a_1 _10760_ (.A1(\sha256cu.msg_scheduler.mreg_11[9] ),
    .A2(_04659_),
    .B1(_04669_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _10761_ (.A(\sha256cu.msg_scheduler.mreg_12[10] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04670_));
 sky130_fd_sc_hd__o211a_1 _10762_ (.A1(\sha256cu.msg_scheduler.mreg_11[10] ),
    .A2(_04659_),
    .B1(_04670_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _10763_ (.A(\sha256cu.msg_scheduler.mreg_12[11] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04671_));
 sky130_fd_sc_hd__o211a_1 _10764_ (.A1(\sha256cu.msg_scheduler.mreg_11[11] ),
    .A2(_04659_),
    .B1(_04671_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00823_));
 sky130_fd_sc_hd__buf_2 _10765_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04672_));
 sky130_fd_sc_hd__or2_1 _10766_ (.A(\sha256cu.msg_scheduler.mreg_12[12] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04673_));
 sky130_fd_sc_hd__o211a_1 _10767_ (.A1(\sha256cu.msg_scheduler.mreg_11[12] ),
    .A2(_04672_),
    .B1(_04673_),
    .C1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _10768_ (.A(\sha256cu.msg_scheduler.mreg_12[13] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04674_));
 sky130_fd_sc_hd__buf_2 _10769_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04675_));
 sky130_fd_sc_hd__o211a_1 _10770_ (.A1(\sha256cu.msg_scheduler.mreg_11[13] ),
    .A2(_04672_),
    .B1(_04674_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00825_));
 sky130_fd_sc_hd__or2_1 _10771_ (.A(\sha256cu.msg_scheduler.mreg_12[14] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04676_));
 sky130_fd_sc_hd__o211a_1 _10772_ (.A1(\sha256cu.msg_scheduler.mreg_11[14] ),
    .A2(_04672_),
    .B1(_04676_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _10773_ (.A(\sha256cu.msg_scheduler.mreg_12[15] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04677_));
 sky130_fd_sc_hd__o211a_1 _10774_ (.A1(\sha256cu.msg_scheduler.mreg_11[15] ),
    .A2(_04672_),
    .B1(_04677_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00827_));
 sky130_fd_sc_hd__or2_1 _10775_ (.A(\sha256cu.msg_scheduler.mreg_12[16] ),
    .B(_04666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04678_));
 sky130_fd_sc_hd__o211a_1 _10776_ (.A1(\sha256cu.msg_scheduler.mreg_11[16] ),
    .A2(_04672_),
    .B1(_04678_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00828_));
 sky130_fd_sc_hd__clkbuf_2 _10777_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04679_));
 sky130_fd_sc_hd__or2_1 _10778_ (.A(\sha256cu.msg_scheduler.mreg_12[17] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04680_));
 sky130_fd_sc_hd__o211a_1 _10779_ (.A1(\sha256cu.msg_scheduler.mreg_11[17] ),
    .A2(_04672_),
    .B1(_04680_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00829_));
 sky130_fd_sc_hd__or2_1 _10780_ (.A(\sha256cu.msg_scheduler.mreg_12[18] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04681_));
 sky130_fd_sc_hd__o211a_1 _10781_ (.A1(\sha256cu.msg_scheduler.mreg_11[18] ),
    .A2(_04672_),
    .B1(_04681_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00830_));
 sky130_fd_sc_hd__or2_1 _10782_ (.A(\sha256cu.msg_scheduler.mreg_12[19] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04682_));
 sky130_fd_sc_hd__o211a_1 _10783_ (.A1(\sha256cu.msg_scheduler.mreg_11[19] ),
    .A2(_04672_),
    .B1(_04682_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _10784_ (.A(\sha256cu.msg_scheduler.mreg_12[20] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04683_));
 sky130_fd_sc_hd__o211a_1 _10785_ (.A1(\sha256cu.msg_scheduler.mreg_11[20] ),
    .A2(_04672_),
    .B1(_04683_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _10786_ (.A(\sha256cu.msg_scheduler.mreg_12[21] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04684_));
 sky130_fd_sc_hd__o211a_1 _10787_ (.A1(\sha256cu.msg_scheduler.mreg_11[21] ),
    .A2(_04672_),
    .B1(_04684_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00833_));
 sky130_fd_sc_hd__clkbuf_4 _10788_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04685_));
 sky130_fd_sc_hd__or2_1 _10789_ (.A(\sha256cu.msg_scheduler.mreg_12[22] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04686_));
 sky130_fd_sc_hd__o211a_1 _10790_ (.A1(\sha256cu.msg_scheduler.mreg_11[22] ),
    .A2(_04685_),
    .B1(_04686_),
    .C1(_04675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00834_));
 sky130_fd_sc_hd__or2_1 _10791_ (.A(\sha256cu.msg_scheduler.mreg_12[23] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_4 _10792_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04688_));
 sky130_fd_sc_hd__o211a_1 _10793_ (.A1(\sha256cu.msg_scheduler.mreg_11[23] ),
    .A2(_04685_),
    .B1(_04687_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00835_));
 sky130_fd_sc_hd__or2_1 _10794_ (.A(\sha256cu.msg_scheduler.mreg_12[24] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04689_));
 sky130_fd_sc_hd__o211a_1 _10795_ (.A1(\sha256cu.msg_scheduler.mreg_11[24] ),
    .A2(_04685_),
    .B1(_04689_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00836_));
 sky130_fd_sc_hd__or2_1 _10796_ (.A(\sha256cu.msg_scheduler.mreg_12[25] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04690_));
 sky130_fd_sc_hd__o211a_1 _10797_ (.A1(\sha256cu.msg_scheduler.mreg_11[25] ),
    .A2(_04685_),
    .B1(_04690_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _10798_ (.A(\sha256cu.msg_scheduler.mreg_12[26] ),
    .B(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04691_));
 sky130_fd_sc_hd__o211a_1 _10799_ (.A1(\sha256cu.msg_scheduler.mreg_11[26] ),
    .A2(_04685_),
    .B1(_04691_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00838_));
 sky130_fd_sc_hd__buf_4 _10800_ (.A(_01566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04692_));
 sky130_fd_sc_hd__or2_1 _10801_ (.A(\sha256cu.msg_scheduler.mreg_12[27] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04693_));
 sky130_fd_sc_hd__o211a_1 _10802_ (.A1(\sha256cu.msg_scheduler.mreg_11[27] ),
    .A2(_04685_),
    .B1(_04693_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00839_));
 sky130_fd_sc_hd__or2_1 _10803_ (.A(\sha256cu.msg_scheduler.mreg_12[28] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04694_));
 sky130_fd_sc_hd__o211a_1 _10804_ (.A1(\sha256cu.msg_scheduler.mreg_11[28] ),
    .A2(_04685_),
    .B1(_04694_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00840_));
 sky130_fd_sc_hd__or2_1 _10805_ (.A(\sha256cu.msg_scheduler.mreg_12[29] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04695_));
 sky130_fd_sc_hd__o211a_1 _10806_ (.A1(\sha256cu.msg_scheduler.mreg_11[29] ),
    .A2(_04685_),
    .B1(_04695_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00841_));
 sky130_fd_sc_hd__or2_1 _10807_ (.A(\sha256cu.msg_scheduler.mreg_12[30] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04696_));
 sky130_fd_sc_hd__o211a_1 _10808_ (.A1(\sha256cu.msg_scheduler.mreg_11[30] ),
    .A2(_04685_),
    .B1(_04696_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _10809_ (.A(\sha256cu.msg_scheduler.mreg_12[31] ),
    .B(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04697_));
 sky130_fd_sc_hd__o211a_1 _10810_ (.A1(\sha256cu.msg_scheduler.mreg_11[31] ),
    .A2(_04685_),
    .B1(_04697_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00843_));
 sky130_fd_sc_hd__clkbuf_4 _10811_ (.A(_01956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04698_));
 sky130_fd_sc_hd__nor2_8 _10812_ (.A(\sha256cu.byte_rdy ),
    .B(_01945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04699_));
 sky130_fd_sc_hd__nand2_2 _10813_ (.A(_04698_),
    .B(_04699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04700_));
 sky130_fd_sc_hd__clkbuf_4 _10814_ (.A(\sha256cu.m_pad_pars.temp_chk ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04701_));
 sky130_fd_sc_hd__clkbuf_4 _10815_ (.A(_04701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04702_));
 sky130_fd_sc_hd__or2_4 _10816_ (.A(\sha256cu.byte_rdy ),
    .B(_01945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04703_));
 sky130_fd_sc_hd__buf_4 _10817_ (.A(_04703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_4 _10818_ (.A(_04704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04705_));
 sky130_fd_sc_hd__nor2_1 _10819_ (.A(_04702_),
    .B(_04705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04706_));
 sky130_fd_sc_hd__or2_1 _10820_ (.A(\sha256cu.m_pad_pars.m_size[3] ),
    .B(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04707_));
 sky130_fd_sc_hd__o211a_1 _10821_ (.A1(_01939_),
    .A2(_04700_),
    .B1(_04707_),
    .C1(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00844_));
 sky130_fd_sc_hd__or2_1 _10822_ (.A(\sha256cu.m_pad_pars.m_size[4] ),
    .B(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_4 _10823_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04709_));
 sky130_fd_sc_hd__o211a_1 _10824_ (.A1(\sha256cu.m_pad_pars.add_512_block[1] ),
    .A2(_04700_),
    .B1(_04708_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00845_));
 sky130_fd_sc_hd__or2_1 _10825_ (.A(\sha256cu.m_pad_pars.m_size[5] ),
    .B(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04710_));
 sky130_fd_sc_hd__o211a_1 _10826_ (.A1(\sha256cu.m_pad_pars.add_512_block[2] ),
    .A2(_04700_),
    .B1(_04710_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00846_));
 sky130_fd_sc_hd__or2_1 _10827_ (.A(\sha256cu.m_pad_pars.m_size[6] ),
    .B(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04711_));
 sky130_fd_sc_hd__o211a_1 _10828_ (.A1(\sha256cu.m_pad_pars.add_512_block[3] ),
    .A2(_04700_),
    .B1(_04711_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00847_));
 sky130_fd_sc_hd__or2_1 _10829_ (.A(\sha256cu.m_pad_pars.m_size[7] ),
    .B(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04712_));
 sky130_fd_sc_hd__o211a_1 _10830_ (.A1(\sha256cu.m_pad_pars.add_512_block[4] ),
    .A2(_04700_),
    .B1(_04712_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00848_));
 sky130_fd_sc_hd__or2_1 _10831_ (.A(\sha256cu.m_pad_pars.m_size[8] ),
    .B(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04713_));
 sky130_fd_sc_hd__o211a_1 _10832_ (.A1(\sha256cu.m_pad_pars.add_512_block[5] ),
    .A2(_04700_),
    .B1(_04713_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00849_));
 sky130_fd_sc_hd__and3_1 _10833_ (.A(\sha256cu.m_pad_pars.m_size[9] ),
    .B(_01994_),
    .C(_04700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04714_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_04714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00850_));
 sky130_fd_sc_hd__a21oi_1 _10835_ (.A1(\sha256cu.msg_scheduler.temp_case ),
    .A2(_04190_),
    .B1(\sha256cu.msg_scheduler.counter_iteration[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04715_));
 sky130_fd_sc_hd__nor2_1 _10836_ (.A(\sha256cu.msg_scheduler.counter_iteration[6] ),
    .B(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04716_));
 sky130_fd_sc_hd__o221ai_1 _10837_ (.A1(_04176_),
    .A2(_04715_),
    .B1(_04716_),
    .B2(\sha256cu.iter_processing.padding_done ),
    .C1(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00851_));
 sky130_fd_sc_hd__a21oi_1 _10838_ (.A1(\sha256cu.msg_scheduler.counter_iteration[6] ),
    .A2(_04185_),
    .B1(_04177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04717_));
 sky130_fd_sc_hd__o21a_1 _10839_ (.A1(\sha256cu.msg_scheduler.counter_iteration[6] ),
    .A2(_04185_),
    .B1(_04717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00852_));
 sky130_fd_sc_hd__and2_1 _10840_ (.A(\sha256cu.m_pad_pars.add_out2[2] ),
    .B(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04718_));
 sky130_fd_sc_hd__o21ai_1 _10841_ (.A1(\sha256cu.m_pad_pars.add_out2[2] ),
    .A2(_01963_),
    .B1(_01966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04719_));
 sky130_fd_sc_hd__nor2_1 _10842_ (.A(_04718_),
    .B(_04719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_1 _10843_ (.A(\sha256cu.m_pad_pars.add_out2[3] ),
    .B(\sha256cu.m_pad_pars.add_out2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04720_));
 sky130_fd_sc_hd__o221a_1 _10844_ (.A1(\sha256cu.m_pad_pars.add_out2[3] ),
    .A2(_04718_),
    .B1(_04720_),
    .B2(_01971_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00854_));
 sky130_fd_sc_hd__clkbuf_2 _10845_ (.A(\sha256cu.m_pad_pars.add_out2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04721_));
 sky130_fd_sc_hd__a31o_1 _10846_ (.A1(\sha256cu.m_pad_pars.add_out2[3] ),
    .A2(\sha256cu.m_pad_pars.add_out2[2] ),
    .A3(_01976_),
    .B1(_04721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04722_));
 sky130_fd_sc_hd__or3b_1 _10847_ (.A(_01980_),
    .B(_04720_),
    .C_N(_04721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04723_));
 sky130_fd_sc_hd__and3_1 _10848_ (.A(_01975_),
    .B(_04722_),
    .C(_04723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04724_));
 sky130_fd_sc_hd__clkbuf_1 _10849_ (.A(_04724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00855_));
 sky130_fd_sc_hd__clkbuf_2 _10850_ (.A(\sha256cu.m_pad_pars.add_out2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04725_));
 sky130_fd_sc_hd__and2b_2 _10851_ (.A_N(\sha256cu.m_pad_pars.add_out2[5] ),
    .B(\sha256cu.m_pad_pars.add_out2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04726_));
 sky130_fd_sc_hd__and3_1 _10852_ (.A(\sha256cu.m_pad_pars.add_out2[3] ),
    .B(\sha256cu.m_pad_pars.add_out2[2] ),
    .C(_04726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04727_));
 sky130_fd_sc_hd__a32o_1 _10853_ (.A1(_04725_),
    .A2(_01966_),
    .A3(_04723_),
    .B1(_04727_),
    .B2(_01987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00856_));
 sky130_fd_sc_hd__and2_1 _10854_ (.A(\sha256cu.m_pad_pars.add_out3[2] ),
    .B(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04728_));
 sky130_fd_sc_hd__o21ai_1 _10855_ (.A1(\sha256cu.m_pad_pars.add_out3[2] ),
    .A2(_01963_),
    .B1(_01966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04729_));
 sky130_fd_sc_hd__nor2_1 _10856_ (.A(_04728_),
    .B(_04729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00857_));
 sky130_fd_sc_hd__nand2_2 _10857_ (.A(\sha256cu.m_pad_pars.add_out3[3] ),
    .B(\sha256cu.m_pad_pars.add_out3[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04730_));
 sky130_fd_sc_hd__o221a_1 _10858_ (.A1(\sha256cu.m_pad_pars.add_out3[3] ),
    .A2(_04728_),
    .B1(_04730_),
    .B2(_01971_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00858_));
 sky130_fd_sc_hd__nor2_1 _10859_ (.A(_01979_),
    .B(_04730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04731_));
 sky130_fd_sc_hd__or2_1 _10860_ (.A(\sha256cu.m_pad_pars.add_out3[4] ),
    .B(_04731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04732_));
 sky130_fd_sc_hd__nand2_1 _10861_ (.A(\sha256cu.m_pad_pars.add_out3[4] ),
    .B(_04731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04733_));
 sky130_fd_sc_hd__and3_1 _10862_ (.A(_01975_),
    .B(_04732_),
    .C(_04733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04734_));
 sky130_fd_sc_hd__clkbuf_1 _10863_ (.A(_04734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00859_));
 sky130_fd_sc_hd__inv_2 _10864_ (.A(\sha256cu.m_pad_pars.add_out3[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04735_));
 sky130_fd_sc_hd__and2_1 _10865_ (.A(\sha256cu.m_pad_pars.add_out3[5] ),
    .B(\sha256cu.m_pad_pars.add_out3[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04736_));
 sky130_fd_sc_hd__and3_1 _10866_ (.A(\sha256cu.m_pad_pars.add_out3[3] ),
    .B(\sha256cu.m_pad_pars.add_out3[2] ),
    .C(_04736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04737_));
 sky130_fd_sc_hd__clkbuf_4 _10867_ (.A(_04737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04738_));
 sky130_fd_sc_hd__and2_1 _10868_ (.A(_01976_),
    .B(_04738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04739_));
 sky130_fd_sc_hd__a211oi_1 _10869_ (.A1(_04735_),
    .A2(_04733_),
    .B1(_04739_),
    .C1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00860_));
 sky130_fd_sc_hd__a31o_1 _10870_ (.A1(\sha256cu.m_pad_pars.add_out3[6] ),
    .A2(_01963_),
    .A3(_04738_),
    .B1(_02002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04740_));
 sky130_fd_sc_hd__o21ba_1 _10871_ (.A1(\sha256cu.m_pad_pars.add_out3[6] ),
    .A2(_04739_),
    .B1_N(_04740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00861_));
 sky130_fd_sc_hd__nor2_1 _10872_ (.A(_02002_),
    .B(_01960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00896_));
 sky130_fd_sc_hd__a22o_1 _10873_ (.A1(\sha256cu.flag_0_15 ),
    .A2(_01966_),
    .B1(_01938_),
    .B2(_00896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00862_));
 sky130_fd_sc_hd__clkbuf_4 _10874_ (.A(_01980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_4 _10875_ (.A(_01987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04742_));
 sky130_fd_sc_hd__inv_2 _10876_ (.A(\sha256cu.m_pad_pars.add_512_block[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_2 _10877_ (.A(_04743_),
    .B(\sha256cu.m_pad_pars.add_512_block[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04744_));
 sky130_fd_sc_hd__or2_1 _10878_ (.A(_04703_),
    .B(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04745_));
 sky130_fd_sc_hd__clkbuf_4 _10879_ (.A(_04745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04746_));
 sky130_fd_sc_hd__buf_4 _10880_ (.A(_04746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04747_));
 sky130_fd_sc_hd__nand2_2 _10881_ (.A(\sha256cu.m_pad_pars.add_512_block[1] ),
    .B(_01939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04748_));
 sky130_fd_sc_hd__or2b_1 _10882_ (.A(\sha256cu.m_pad_pars.add_512_block[2] ),
    .B_N(\sha256cu.m_pad_pars.add_512_block[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04749_));
 sky130_fd_sc_hd__or2_1 _10883_ (.A(_04748_),
    .B(_04749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04750_));
 sky130_fd_sc_hd__buf_2 _10884_ (.A(_04750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04751_));
 sky130_fd_sc_hd__or2b_1 _10885_ (.A(_01939_),
    .B_N(\sha256cu.m_pad_pars.add_512_block[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04752_));
 sky130_fd_sc_hd__or2_2 _10886_ (.A(_04749_),
    .B(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04753_));
 sky130_fd_sc_hd__o21a_1 _10887_ (.A1(_04702_),
    .A2(_04751_),
    .B1(_04753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04754_));
 sky130_fd_sc_hd__and2b_1 _10888_ (.A_N(\sha256cu.m_pad_pars.add_out3[2] ),
    .B(\sha256cu.m_pad_pars.add_out3[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04755_));
 sky130_fd_sc_hd__and2_2 _10889_ (.A(_04735_),
    .B(\sha256cu.m_pad_pars.add_out3[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04756_));
 sky130_fd_sc_hd__o211a_2 _10890_ (.A1(_04747_),
    .A2(_04754_),
    .B1(_04755_),
    .C1(_04756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04757_));
 sky130_fd_sc_hd__or2_2 _10891_ (.A(_01940_),
    .B(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04758_));
 sky130_fd_sc_hd__or2_2 _10892_ (.A(_04704_),
    .B(_04758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04759_));
 sky130_fd_sc_hd__nor2_2 _10893_ (.A(_04748_),
    .B(_01940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_2 _10894_ (.A(_04699_),
    .B(_04760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04761_));
 sky130_fd_sc_hd__nor2_1 _10895_ (.A(_01943_),
    .B(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04762_));
 sky130_fd_sc_hd__a2bb2o_1 _10896_ (.A1_N(_01943_),
    .A2_N(_04759_),
    .B1(_04762_),
    .B2(_04698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04763_));
 sky130_fd_sc_hd__nor2_2 _10897_ (.A(\sha256cu.m_pad_pars.add_out3[3] ),
    .B(\sha256cu.m_pad_pars.add_out3[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04764_));
 sky130_fd_sc_hd__and4bb_4 _10898_ (.A_N(_04763_),
    .B_N(\sha256cu.m_pad_pars.add_out3[4] ),
    .C(_04735_),
    .D(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04765_));
 sky130_fd_sc_hd__nor2_1 _10899_ (.A(\sha256cu.m_pad_pars.add_out3[5] ),
    .B(\sha256cu.m_pad_pars.add_out3[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04766_));
 sky130_fd_sc_hd__and2b_1 _10900_ (.A_N(\sha256cu.m_pad_pars.add_out3[3] ),
    .B(\sha256cu.m_pad_pars.add_out3[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04767_));
 sky130_fd_sc_hd__nand2_4 _10901_ (.A(_01944_),
    .B(_04699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04768_));
 sky130_fd_sc_hd__buf_4 _10902_ (.A(_04768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04769_));
 sky130_fd_sc_hd__or2_2 _10903_ (.A(_04748_),
    .B(_01953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04770_));
 sky130_fd_sc_hd__or2_2 _10904_ (.A(_01953_),
    .B(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04771_));
 sky130_fd_sc_hd__or2_1 _10905_ (.A(_04768_),
    .B(_04771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04772_));
 sky130_fd_sc_hd__o31a_1 _10906_ (.A1(_04702_),
    .A2(_04769_),
    .A3(_04770_),
    .B1(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04773_));
 sky130_fd_sc_hd__and3_2 _10907_ (.A(_04766_),
    .B(_04767_),
    .C(_04773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04774_));
 sky130_fd_sc_hd__nor2_2 _10908_ (.A(_04701_),
    .B(_04768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04775_));
 sky130_fd_sc_hd__nand2_2 _10909_ (.A(\sha256cu.m_pad_pars.add_512_block[3] ),
    .B(\sha256cu.m_pad_pars.add_512_block[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04776_));
 sky130_fd_sc_hd__nor2_2 _10910_ (.A(_04748_),
    .B(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04777_));
 sky130_fd_sc_hd__nand2_1 _10911_ (.A(_04775_),
    .B(_04777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04778_));
 sky130_fd_sc_hd__or2_2 _10912_ (.A(_04752_),
    .B(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04779_));
 sky130_fd_sc_hd__or2_1 _10913_ (.A(_04768_),
    .B(_04779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04780_));
 sky130_fd_sc_hd__and4b_2 _10914_ (.A_N(_04730_),
    .B(_04766_),
    .C(_04778_),
    .D(_04780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04781_));
 sky130_fd_sc_hd__a22o_1 _10915_ (.A1(\sha256cu.m_pad_pars.block_512[7][0] ),
    .A2(_04774_),
    .B1(_04781_),
    .B2(\sha256cu.m_pad_pars.block_512[15][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04782_));
 sky130_fd_sc_hd__a221o_1 _10916_ (.A1(\sha256cu.m_pad_pars.block_512[27][0] ),
    .A2(_04757_),
    .B1(_04765_),
    .B2(\sha256cu.m_pad_pars.block_512[3][0] ),
    .C1(_04782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04783_));
 sky130_fd_sc_hd__nand2_1 _10917_ (.A(_04755_),
    .B(_04766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04784_));
 sky130_fd_sc_hd__nor2_2 _10918_ (.A(_04749_),
    .B(_04752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04785_));
 sky130_fd_sc_hd__nor2_4 _10919_ (.A(_01943_),
    .B(_04703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2_4 _10920_ (.A(_01956_),
    .B(_04786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04787_));
 sky130_fd_sc_hd__nor2_1 _10921_ (.A(_04751_),
    .B(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04788_));
 sky130_fd_sc_hd__a21o_1 _10922_ (.A1(_04785_),
    .A2(_04786_),
    .B1(_04788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04789_));
 sky130_fd_sc_hd__nor2_4 _10923_ (.A(_04784_),
    .B(_04789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04790_));
 sky130_fd_sc_hd__or2_4 _10924_ (.A(_04743_),
    .B(\sha256cu.m_pad_pars.add_512_block[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04791_));
 sky130_fd_sc_hd__or2_2 _10925_ (.A(\sha256cu.m_pad_pars.temp_chk ),
    .B(_04791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04792_));
 sky130_fd_sc_hd__or2_1 _10926_ (.A(_04703_),
    .B(_04792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04793_));
 sky130_fd_sc_hd__buf_2 _10927_ (.A(_04793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04794_));
 sky130_fd_sc_hd__nor2_2 _10928_ (.A(_04770_),
    .B(_04794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04795_));
 sky130_fd_sc_hd__or2_1 _10929_ (.A(_04703_),
    .B(_04771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04796_));
 sky130_fd_sc_hd__or2_1 _10930_ (.A(_04796_),
    .B(_04791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04797_));
 sky130_fd_sc_hd__nor2_1 _10931_ (.A(_04735_),
    .B(\sha256cu.m_pad_pars.add_out3[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04798_));
 sky130_fd_sc_hd__and2_1 _10932_ (.A(_04767_),
    .B(_04798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04799_));
 sky130_fd_sc_hd__and3b_2 _10933_ (.A_N(_04795_),
    .B(_04797_),
    .C(_04799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04800_));
 sky130_fd_sc_hd__nor2_4 _10934_ (.A(_04704_),
    .B(_04791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _10935_ (.A(_04751_),
    .B(_04794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04802_));
 sky130_fd_sc_hd__a21oi_1 _10936_ (.A1(_04785_),
    .A2(_04801_),
    .B1(_04802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04803_));
 sky130_fd_sc_hd__and3_2 _10937_ (.A(_04755_),
    .B(_04798_),
    .C(_04803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04804_));
 sky130_fd_sc_hd__or2_1 _10938_ (.A(\sha256cu.m_pad_pars.add_512_block[6] ),
    .B(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04805_));
 sky130_fd_sc_hd__or2_1 _10939_ (.A(\sha256cu.m_pad_pars.temp_chk ),
    .B(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04806_));
 sky130_fd_sc_hd__clkbuf_4 _10940_ (.A(_04806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04807_));
 sky130_fd_sc_hd__or2_2 _10941_ (.A(_04748_),
    .B(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04808_));
 sky130_fd_sc_hd__o22a_1 _10942_ (.A1(_04805_),
    .A2(_04779_),
    .B1(_04807_),
    .B2(_04808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04809_));
 sky130_fd_sc_hd__and3_1 _10943_ (.A(\sha256cu.m_pad_pars.add_out3[3] ),
    .B(\sha256cu.m_pad_pars.add_out3[2] ),
    .C(_04756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04810_));
 sky130_fd_sc_hd__o21a_2 _10944_ (.A1(_04704_),
    .A2(_04809_),
    .B1(_04810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04811_));
 sky130_fd_sc_hd__a22o_1 _10945_ (.A1(\sha256cu.m_pad_pars.block_512[43][0] ),
    .A2(_04804_),
    .B1(_04811_),
    .B2(\sha256cu.m_pad_pars.block_512[31][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04812_));
 sky130_fd_sc_hd__a221o_1 _10946_ (.A1(\sha256cu.m_pad_pars.block_512[11][0] ),
    .A2(_04790_),
    .B1(_04800_),
    .B2(\sha256cu.m_pad_pars.block_512[39][0] ),
    .C1(_04812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04813_));
 sky130_fd_sc_hd__or2_1 _10947_ (.A(_04735_),
    .B(\sha256cu.m_pad_pars.add_out3[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04814_));
 sky130_fd_sc_hd__or2_1 _10948_ (.A(_04748_),
    .B(_01940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04815_));
 sky130_fd_sc_hd__nor2_1 _10949_ (.A(_04815_),
    .B(_04794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04816_));
 sky130_fd_sc_hd__o21bai_2 _10950_ (.A1(_04759_),
    .A2(_04791_),
    .B1_N(_04816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04817_));
 sky130_fd_sc_hd__nor4_4 _10951_ (.A(\sha256cu.m_pad_pars.add_out3[3] ),
    .B(\sha256cu.m_pad_pars.add_out3[2] ),
    .C(_04814_),
    .D(_04817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04818_));
 sky130_fd_sc_hd__or2_2 _10952_ (.A(\sha256cu.m_pad_pars.add_512_block[6] ),
    .B(_04791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04819_));
 sky130_fd_sc_hd__o22a_1 _10953_ (.A1(_04779_),
    .A2(_04819_),
    .B1(_04792_),
    .B2(_04808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04820_));
 sky130_fd_sc_hd__nor2_1 _10954_ (.A(_04730_),
    .B(_04814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04821_));
 sky130_fd_sc_hd__o21a_2 _10955_ (.A1(_04705_),
    .A2(_04820_),
    .B1(_04821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04822_));
 sky130_fd_sc_hd__nor2_2 _10956_ (.A(_01952_),
    .B(_04759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_4 _10957_ (.A(_01956_),
    .B(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04824_));
 sky130_fd_sc_hd__nor2_2 _10958_ (.A(_04761_),
    .B(_04824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04825_));
 sky130_fd_sc_hd__and4bb_4 _10959_ (.A_N(_04823_),
    .B_N(_04825_),
    .C(_04736_),
    .D(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04826_));
 sky130_fd_sc_hd__o32a_1 _10960_ (.A1(_04705_),
    .A2(_04770_),
    .A3(_04807_),
    .B1(_04746_),
    .B2(_04771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04827_));
 sky130_fd_sc_hd__and3_2 _10961_ (.A(_04756_),
    .B(_04767_),
    .C(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04828_));
 sky130_fd_sc_hd__and3_2 _10962_ (.A(_01919_),
    .B(_04736_),
    .C(_04755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04829_));
 sky130_fd_sc_hd__o22a_1 _10963_ (.A1(_04746_),
    .A2(_04758_),
    .B1(_04761_),
    .B2(_04807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04830_));
 sky130_fd_sc_hd__and3_2 _10964_ (.A(_04756_),
    .B(_04764_),
    .C(_04830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04831_));
 sky130_fd_sc_hd__or3_1 _10965_ (.A(_01917_),
    .B(_01951_),
    .C(_04771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04832_));
 sky130_fd_sc_hd__and3_2 _10966_ (.A(_04736_),
    .B(_04767_),
    .C(_04832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04833_));
 sky130_fd_sc_hd__a32o_1 _10967_ (.A1(\sha256cu.m_pad_pars.block_512[63][0] ),
    .A2(_01919_),
    .A3(_04738_),
    .B1(_04833_),
    .B2(\sha256cu.m_pad_pars.block_512[55][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04834_));
 sky130_fd_sc_hd__a221o_1 _10968_ (.A1(\sha256cu.m_pad_pars.block_512[59][0] ),
    .A2(_04829_),
    .B1(_04831_),
    .B2(\sha256cu.m_pad_pars.block_512[19][0] ),
    .C1(_04834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04835_));
 sky130_fd_sc_hd__a221o_1 _10969_ (.A1(\sha256cu.m_pad_pars.block_512[51][0] ),
    .A2(_04826_),
    .B1(_04828_),
    .B2(\sha256cu.m_pad_pars.block_512[23][0] ),
    .C1(_04835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04836_));
 sky130_fd_sc_hd__a221o_1 _10970_ (.A1(\sha256cu.m_pad_pars.block_512[35][0] ),
    .A2(_04818_),
    .B1(_04822_),
    .B2(\sha256cu.m_pad_pars.block_512[47][0] ),
    .C1(_04836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04837_));
 sky130_fd_sc_hd__or2_1 _10971_ (.A(_04813_),
    .B(_04837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04838_));
 sky130_fd_sc_hd__or2_1 _10972_ (.A(_04783_),
    .B(_04838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04839_));
 sky130_fd_sc_hd__a22o_1 _10973_ (.A1(\sha256cu.data_in_padd[0] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_04839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00863_));
 sky130_fd_sc_hd__buf_4 _10974_ (.A(_01963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04840_));
 sky130_fd_sc_hd__a22o_1 _10975_ (.A1(\sha256cu.m_pad_pars.block_512[7][1] ),
    .A2(_04774_),
    .B1(_04781_),
    .B2(\sha256cu.m_pad_pars.block_512[15][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04841_));
 sky130_fd_sc_hd__a211o_1 _10976_ (.A1(\sha256cu.m_pad_pars.block_512[3][1] ),
    .A2(_04765_),
    .B1(_04841_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04842_));
 sky130_fd_sc_hd__a32o_1 _10977_ (.A1(\sha256cu.m_pad_pars.block_512[63][1] ),
    .A2(_01920_),
    .A3(_04738_),
    .B1(_04833_),
    .B2(\sha256cu.m_pad_pars.block_512[55][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04843_));
 sky130_fd_sc_hd__a221o_1 _10978_ (.A1(\sha256cu.m_pad_pars.block_512[11][1] ),
    .A2(_04790_),
    .B1(_04831_),
    .B2(\sha256cu.m_pad_pars.block_512[19][1] ),
    .C1(_04843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04844_));
 sky130_fd_sc_hd__a221o_1 _10979_ (.A1(\sha256cu.m_pad_pars.block_512[27][1] ),
    .A2(_04757_),
    .B1(_04828_),
    .B2(\sha256cu.m_pad_pars.block_512[23][1] ),
    .C1(_04844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04845_));
 sky130_fd_sc_hd__a22o_1 _10980_ (.A1(\sha256cu.m_pad_pars.block_512[39][1] ),
    .A2(_04800_),
    .B1(_04826_),
    .B2(\sha256cu.m_pad_pars.block_512[51][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04846_));
 sky130_fd_sc_hd__a22o_1 _10981_ (.A1(\sha256cu.m_pad_pars.block_512[59][1] ),
    .A2(_04829_),
    .B1(_04822_),
    .B2(\sha256cu.m_pad_pars.block_512[47][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04847_));
 sky130_fd_sc_hd__a21o_1 _10982_ (.A1(\sha256cu.m_pad_pars.block_512[43][1] ),
    .A2(_04804_),
    .B1(_04847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04848_));
 sky130_fd_sc_hd__a211o_1 _10983_ (.A1(\sha256cu.m_pad_pars.block_512[35][1] ),
    .A2(_04818_),
    .B1(_04846_),
    .C1(_04848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04849_));
 sky130_fd_sc_hd__a211o_1 _10984_ (.A1(\sha256cu.m_pad_pars.block_512[31][1] ),
    .A2(_04811_),
    .B1(_04845_),
    .C1(_04849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04850_));
 sky130_fd_sc_hd__o221a_1 _10985_ (.A1(\sha256cu.data_in_padd[1] ),
    .A2(_04840_),
    .B1(_04842_),
    .B2(_04850_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00864_));
 sky130_fd_sc_hd__a22o_1 _10986_ (.A1(\sha256cu.m_pad_pars.block_512[3][2] ),
    .A2(_04765_),
    .B1(_04774_),
    .B2(\sha256cu.m_pad_pars.block_512[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04851_));
 sky130_fd_sc_hd__a211o_1 _10987_ (.A1(\sha256cu.m_pad_pars.block_512[15][2] ),
    .A2(_04781_),
    .B1(_04851_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04852_));
 sky130_fd_sc_hd__a22o_1 _10988_ (.A1(\sha256cu.m_pad_pars.block_512[31][2] ),
    .A2(_04811_),
    .B1(_04822_),
    .B2(\sha256cu.m_pad_pars.block_512[47][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04853_));
 sky130_fd_sc_hd__and2_1 _10989_ (.A(\sha256cu.m_pad_pars.block_512[59][2] ),
    .B(_04829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04854_));
 sky130_fd_sc_hd__a221o_1 _10990_ (.A1(\sha256cu.m_pad_pars.block_512[39][2] ),
    .A2(_04800_),
    .B1(_04831_),
    .B2(\sha256cu.m_pad_pars.block_512[19][2] ),
    .C1(_04854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04855_));
 sky130_fd_sc_hd__a32o_1 _10991_ (.A1(\sha256cu.m_pad_pars.block_512[63][2] ),
    .A2(_01920_),
    .A3(_04738_),
    .B1(_04833_),
    .B2(\sha256cu.m_pad_pars.block_512[55][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04856_));
 sky130_fd_sc_hd__a221o_1 _10992_ (.A1(\sha256cu.m_pad_pars.block_512[27][2] ),
    .A2(_04757_),
    .B1(_04790_),
    .B2(\sha256cu.m_pad_pars.block_512[11][2] ),
    .C1(_04856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04857_));
 sky130_fd_sc_hd__a221o_1 _10993_ (.A1(\sha256cu.m_pad_pars.block_512[43][2] ),
    .A2(_04804_),
    .B1(_04828_),
    .B2(\sha256cu.m_pad_pars.block_512[23][2] ),
    .C1(_04857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04858_));
 sky130_fd_sc_hd__a211o_1 _10994_ (.A1(\sha256cu.m_pad_pars.block_512[35][2] ),
    .A2(_04818_),
    .B1(_04855_),
    .C1(_04858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04859_));
 sky130_fd_sc_hd__a211o_1 _10995_ (.A1(\sha256cu.m_pad_pars.block_512[51][2] ),
    .A2(_04826_),
    .B1(_04853_),
    .C1(_04859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04860_));
 sky130_fd_sc_hd__o221a_1 _10996_ (.A1(\sha256cu.data_in_padd[2] ),
    .A2(_04840_),
    .B1(_04852_),
    .B2(_04860_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\sha256cu.m_pad_pars.m_size[3] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][3] ),
    .S(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04861_));
 sky130_fd_sc_hd__a22o_1 _10998_ (.A1(\sha256cu.m_pad_pars.block_512[59][3] ),
    .A2(_04829_),
    .B1(_04833_),
    .B2(\sha256cu.m_pad_pars.block_512[55][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04862_));
 sky130_fd_sc_hd__a221o_1 _10999_ (.A1(\sha256cu.m_pad_pars.block_512[31][3] ),
    .A2(_04811_),
    .B1(_04861_),
    .B2(_04738_),
    .C1(_04862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04863_));
 sky130_fd_sc_hd__a221o_1 _11000_ (.A1(\sha256cu.m_pad_pars.block_512[51][3] ),
    .A2(_04826_),
    .B1(_04822_),
    .B2(\sha256cu.m_pad_pars.block_512[47][3] ),
    .C1(_04863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04864_));
 sky130_fd_sc_hd__a221o_1 _11001_ (.A1(\sha256cu.m_pad_pars.block_512[27][3] ),
    .A2(_04757_),
    .B1(_04804_),
    .B2(\sha256cu.m_pad_pars.block_512[43][3] ),
    .C1(_04864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04865_));
 sky130_fd_sc_hd__a22o_1 _11002_ (.A1(\sha256cu.m_pad_pars.block_512[3][3] ),
    .A2(_04765_),
    .B1(_04774_),
    .B2(\sha256cu.m_pad_pars.block_512[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04866_));
 sky130_fd_sc_hd__a221o_1 _11003_ (.A1(\sha256cu.m_pad_pars.block_512[23][3] ),
    .A2(_04828_),
    .B1(_04818_),
    .B2(\sha256cu.m_pad_pars.block_512[35][3] ),
    .C1(_04866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04867_));
 sky130_fd_sc_hd__a22o_1 _11004_ (.A1(\sha256cu.m_pad_pars.block_512[11][3] ),
    .A2(_04790_),
    .B1(_04831_),
    .B2(\sha256cu.m_pad_pars.block_512[19][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04868_));
 sky130_fd_sc_hd__a22o_1 _11005_ (.A1(\sha256cu.m_pad_pars.block_512[15][3] ),
    .A2(_04781_),
    .B1(_04800_),
    .B2(\sha256cu.m_pad_pars.block_512[39][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04869_));
 sky130_fd_sc_hd__or4_2 _11006_ (.A(_04865_),
    .B(_04867_),
    .C(_04868_),
    .D(_04869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04870_));
 sky130_fd_sc_hd__or2_1 _11007_ (.A(\sha256cu.data_in_padd[3] ),
    .B(_01963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04871_));
 sky130_fd_sc_hd__o211a_1 _11008_ (.A1(_01971_),
    .A2(_04870_),
    .B1(_04871_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(\sha256cu.m_pad_pars.m_size[4] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][4] ),
    .S(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04872_));
 sky130_fd_sc_hd__a22o_1 _11010_ (.A1(\sha256cu.m_pad_pars.block_512[59][4] ),
    .A2(_04829_),
    .B1(_04833_),
    .B2(\sha256cu.m_pad_pars.block_512[55][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04873_));
 sky130_fd_sc_hd__a221o_1 _11011_ (.A1(\sha256cu.m_pad_pars.block_512[31][4] ),
    .A2(_04811_),
    .B1(_04872_),
    .B2(_04738_),
    .C1(_04873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04874_));
 sky130_fd_sc_hd__a221o_1 _11012_ (.A1(\sha256cu.m_pad_pars.block_512[51][4] ),
    .A2(_04826_),
    .B1(_04822_),
    .B2(\sha256cu.m_pad_pars.block_512[47][4] ),
    .C1(_04874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04875_));
 sky130_fd_sc_hd__a221o_1 _11013_ (.A1(\sha256cu.m_pad_pars.block_512[27][4] ),
    .A2(_04757_),
    .B1(_04804_),
    .B2(\sha256cu.m_pad_pars.block_512[43][4] ),
    .C1(_04875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04876_));
 sky130_fd_sc_hd__a22o_1 _11014_ (.A1(\sha256cu.m_pad_pars.block_512[3][4] ),
    .A2(_04765_),
    .B1(_04774_),
    .B2(\sha256cu.m_pad_pars.block_512[7][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04877_));
 sky130_fd_sc_hd__a221o_1 _11015_ (.A1(\sha256cu.m_pad_pars.block_512[23][4] ),
    .A2(_04828_),
    .B1(_04818_),
    .B2(\sha256cu.m_pad_pars.block_512[35][4] ),
    .C1(_04877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04878_));
 sky130_fd_sc_hd__a22o_1 _11016_ (.A1(\sha256cu.m_pad_pars.block_512[11][4] ),
    .A2(_04790_),
    .B1(_04831_),
    .B2(\sha256cu.m_pad_pars.block_512[19][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04879_));
 sky130_fd_sc_hd__a22o_1 _11017_ (.A1(\sha256cu.m_pad_pars.block_512[15][4] ),
    .A2(_04781_),
    .B1(_04800_),
    .B2(\sha256cu.m_pad_pars.block_512[39][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04880_));
 sky130_fd_sc_hd__or4_2 _11018_ (.A(_04876_),
    .B(_04878_),
    .C(_04879_),
    .D(_04880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04881_));
 sky130_fd_sc_hd__or2_1 _11019_ (.A(\sha256cu.data_in_padd[4] ),
    .B(_01963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04882_));
 sky130_fd_sc_hd__o211a_1 _11020_ (.A1(_01971_),
    .A2(_04881_),
    .B1(_04882_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(\sha256cu.m_pad_pars.m_size[5] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][5] ),
    .S(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04883_));
 sky130_fd_sc_hd__a22o_1 _11022_ (.A1(\sha256cu.m_pad_pars.block_512[31][5] ),
    .A2(_04811_),
    .B1(_04883_),
    .B2(_04738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04884_));
 sky130_fd_sc_hd__a221o_1 _11023_ (.A1(\sha256cu.m_pad_pars.block_512[59][5] ),
    .A2(_04829_),
    .B1(_04833_),
    .B2(\sha256cu.m_pad_pars.block_512[55][5] ),
    .C1(_04884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04885_));
 sky130_fd_sc_hd__a221o_1 _11024_ (.A1(\sha256cu.m_pad_pars.block_512[51][5] ),
    .A2(_04826_),
    .B1(_04822_),
    .B2(\sha256cu.m_pad_pars.block_512[47][5] ),
    .C1(_04885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04886_));
 sky130_fd_sc_hd__a221o_1 _11025_ (.A1(\sha256cu.m_pad_pars.block_512[27][5] ),
    .A2(_04757_),
    .B1(_04804_),
    .B2(\sha256cu.m_pad_pars.block_512[43][5] ),
    .C1(_04886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04887_));
 sky130_fd_sc_hd__a22o_1 _11026_ (.A1(\sha256cu.m_pad_pars.block_512[3][5] ),
    .A2(_04765_),
    .B1(_04774_),
    .B2(\sha256cu.m_pad_pars.block_512[7][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04888_));
 sky130_fd_sc_hd__a221o_1 _11027_ (.A1(\sha256cu.m_pad_pars.block_512[23][5] ),
    .A2(_04828_),
    .B1(_04818_),
    .B2(\sha256cu.m_pad_pars.block_512[35][5] ),
    .C1(_04888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04889_));
 sky130_fd_sc_hd__a22o_1 _11028_ (.A1(\sha256cu.m_pad_pars.block_512[11][5] ),
    .A2(_04790_),
    .B1(_04831_),
    .B2(\sha256cu.m_pad_pars.block_512[19][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04890_));
 sky130_fd_sc_hd__a22o_1 _11029_ (.A1(\sha256cu.m_pad_pars.block_512[15][5] ),
    .A2(_04781_),
    .B1(_04800_),
    .B2(\sha256cu.m_pad_pars.block_512[39][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04891_));
 sky130_fd_sc_hd__or4_2 _11030_ (.A(_04887_),
    .B(_04889_),
    .C(_04890_),
    .D(_04891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04892_));
 sky130_fd_sc_hd__or2_1 _11031_ (.A(\sha256cu.data_in_padd[5] ),
    .B(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04893_));
 sky130_fd_sc_hd__o211a_1 _11032_ (.A1(_01971_),
    .A2(_04892_),
    .B1(_04893_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(\sha256cu.m_pad_pars.m_size[6] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][6] ),
    .S(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04894_));
 sky130_fd_sc_hd__a22o_1 _11034_ (.A1(\sha256cu.m_pad_pars.block_512[35][6] ),
    .A2(_04818_),
    .B1(_04894_),
    .B2(_04738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04895_));
 sky130_fd_sc_hd__a221o_1 _11035_ (.A1(\sha256cu.m_pad_pars.block_512[59][6] ),
    .A2(_04829_),
    .B1(_04833_),
    .B2(\sha256cu.m_pad_pars.block_512[55][6] ),
    .C1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04896_));
 sky130_fd_sc_hd__a221o_1 _11036_ (.A1(\sha256cu.m_pad_pars.block_512[15][6] ),
    .A2(_04781_),
    .B1(_04790_),
    .B2(\sha256cu.m_pad_pars.block_512[11][6] ),
    .C1(_04896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04897_));
 sky130_fd_sc_hd__a22o_1 _11037_ (.A1(\sha256cu.m_pad_pars.block_512[27][6] ),
    .A2(_04757_),
    .B1(_04804_),
    .B2(\sha256cu.m_pad_pars.block_512[43][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04898_));
 sky130_fd_sc_hd__a22o_1 _11038_ (.A1(\sha256cu.m_pad_pars.block_512[31][6] ),
    .A2(_04811_),
    .B1(_04828_),
    .B2(\sha256cu.m_pad_pars.block_512[23][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04899_));
 sky130_fd_sc_hd__a221o_1 _11039_ (.A1(\sha256cu.m_pad_pars.block_512[39][6] ),
    .A2(_04800_),
    .B1(_04831_),
    .B2(\sha256cu.m_pad_pars.block_512[19][6] ),
    .C1(_04899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04900_));
 sky130_fd_sc_hd__a22o_1 _11040_ (.A1(\sha256cu.m_pad_pars.block_512[7][6] ),
    .A2(_04774_),
    .B1(_04822_),
    .B2(\sha256cu.m_pad_pars.block_512[47][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04901_));
 sky130_fd_sc_hd__a221o_1 _11041_ (.A1(\sha256cu.m_pad_pars.block_512[3][6] ),
    .A2(_04765_),
    .B1(_04826_),
    .B2(\sha256cu.m_pad_pars.block_512[51][6] ),
    .C1(_04901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04902_));
 sky130_fd_sc_hd__or4_2 _11042_ (.A(_04897_),
    .B(_04898_),
    .C(_04900_),
    .D(_04902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04903_));
 sky130_fd_sc_hd__or2_1 _11043_ (.A(\sha256cu.data_in_padd[6] ),
    .B(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04904_));
 sky130_fd_sc_hd__o211a_1 _11044_ (.A1(_01971_),
    .A2(_04903_),
    .B1(_04904_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(\sha256cu.m_pad_pars.m_size[7] ),
    .A1(\sha256cu.m_pad_pars.block_512[63][7] ),
    .S(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04905_));
 sky130_fd_sc_hd__a22o_1 _11046_ (.A1(\sha256cu.m_pad_pars.block_512[55][7] ),
    .A2(_04833_),
    .B1(_04905_),
    .B2(_04738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04906_));
 sky130_fd_sc_hd__clkbuf_4 _11047_ (.A(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04907_));
 sky130_fd_sc_hd__nor2_4 _11048_ (.A(_04704_),
    .B(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04908_));
 sky130_fd_sc_hd__nand2_1 _11049_ (.A(_04908_),
    .B(_04777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04909_));
 sky130_fd_sc_hd__nor2_1 _11050_ (.A(_04702_),
    .B(_04909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04910_));
 sky130_fd_sc_hd__o22a_1 _11051_ (.A1(_04907_),
    .A2(_04779_),
    .B1(_04910_),
    .B2(\sha256cu.m_pad_pars.block_512[31][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04911_));
 sky130_fd_sc_hd__or2_4 _11052_ (.A(_04704_),
    .B(_04791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04912_));
 sky130_fd_sc_hd__buf_4 _11053_ (.A(_04912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04913_));
 sky130_fd_sc_hd__o22a_1 _11054_ (.A1(_04753_),
    .A2(_04913_),
    .B1(_04802_),
    .B2(\sha256cu.m_pad_pars.block_512[43][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04914_));
 sky130_fd_sc_hd__and3_1 _11055_ (.A(_04755_),
    .B(_04798_),
    .C(_04914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04915_));
 sky130_fd_sc_hd__a21o_1 _11056_ (.A1(_04810_),
    .A2(_04911_),
    .B1(_04915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04916_));
 sky130_fd_sc_hd__buf_4 _11057_ (.A(_04913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04917_));
 sky130_fd_sc_hd__nor2_1 _11058_ (.A(_04808_),
    .B(_04794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04918_));
 sky130_fd_sc_hd__o22a_1 _11059_ (.A1(_04779_),
    .A2(_04917_),
    .B1(_04918_),
    .B2(\sha256cu.m_pad_pars.block_512[47][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04919_));
 sky130_fd_sc_hd__o22a_1 _11060_ (.A1(_04758_),
    .A2(_04913_),
    .B1(_04816_),
    .B2(\sha256cu.m_pad_pars.block_512[35][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04920_));
 sky130_fd_sc_hd__and3_1 _11061_ (.A(_04764_),
    .B(_04798_),
    .C(_04920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04921_));
 sky130_fd_sc_hd__nor2_1 _11062_ (.A(_04770_),
    .B(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04922_));
 sky130_fd_sc_hd__o21a_1 _11063_ (.A1(\sha256cu.m_pad_pars.block_512[7][7] ),
    .A2(_04922_),
    .B1(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04923_));
 sky130_fd_sc_hd__nor2_1 _11064_ (.A(_04748_),
    .B(_01953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04924_));
 sky130_fd_sc_hd__nor2_1 _11065_ (.A(_04701_),
    .B(_04744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04925_));
 sky130_fd_sc_hd__a31o_1 _11066_ (.A1(_04699_),
    .A2(_04924_),
    .A3(_04925_),
    .B1(\sha256cu.m_pad_pars.block_512[23][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04926_));
 sky130_fd_sc_hd__o21a_1 _11067_ (.A1(_04747_),
    .A2(_04771_),
    .B1(_04926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04927_));
 sky130_fd_sc_hd__and3_1 _11068_ (.A(_04756_),
    .B(_04767_),
    .C(_04927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04928_));
 sky130_fd_sc_hd__a31o_1 _11069_ (.A1(_04766_),
    .A2(_04767_),
    .A3(_04923_),
    .B1(_04928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04929_));
 sky130_fd_sc_hd__a211o_1 _11070_ (.A1(_04821_),
    .A2(_04919_),
    .B1(_04921_),
    .C1(_04929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04930_));
 sky130_fd_sc_hd__a2111o_1 _11071_ (.A1(\sha256cu.m_pad_pars.block_512[59][7] ),
    .A2(_04829_),
    .B1(_04906_),
    .C1(_04916_),
    .D1(_04930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04931_));
 sky130_fd_sc_hd__o21ba_1 _11072_ (.A1(\sha256cu.m_pad_pars.block_512[51][7] ),
    .A2(_04825_),
    .B1_N(_04823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04932_));
 sky130_fd_sc_hd__buf_4 _11073_ (.A(_04769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04933_));
 sky130_fd_sc_hd__a21oi_1 _11074_ (.A1(_04760_),
    .A2(_04775_),
    .B1(\sha256cu.m_pad_pars.block_512[3][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04934_));
 sky130_fd_sc_hd__o21ba_1 _11075_ (.A1(_04758_),
    .A2(_04933_),
    .B1_N(_04934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04935_));
 sky130_fd_sc_hd__o21a_1 _11076_ (.A1(\sha256cu.m_pad_pars.block_512[39][7] ),
    .A2(_04795_),
    .B1(_04797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04936_));
 sky130_fd_sc_hd__inv_2 _11077_ (.A(\sha256cu.m_pad_pars.block_512[15][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04937_));
 sky130_fd_sc_hd__a21bo_1 _11078_ (.A1(_04937_),
    .A2(_04778_),
    .B1_N(_04780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04938_));
 sky130_fd_sc_hd__or4_1 _11079_ (.A(\sha256cu.m_pad_pars.add_out3[5] ),
    .B(\sha256cu.m_pad_pars.add_out3[4] ),
    .C(_04730_),
    .D(_04938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04939_));
 sky130_fd_sc_hd__a21bo_1 _11080_ (.A1(_04799_),
    .A2(_04936_),
    .B1_N(_04939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04940_));
 sky130_fd_sc_hd__a311o_1 _11081_ (.A1(_04764_),
    .A2(_04766_),
    .A3(_04935_),
    .B1(_04940_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04941_));
 sky130_fd_sc_hd__nor2_1 _11082_ (.A(_04761_),
    .B(_04807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04942_));
 sky130_fd_sc_hd__o22a_1 _11083_ (.A1(_04907_),
    .A2(_04758_),
    .B1(_04942_),
    .B2(\sha256cu.m_pad_pars.block_512[19][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04943_));
 sky130_fd_sc_hd__and3b_1 _11084_ (.A_N(_04751_),
    .B(_04698_),
    .C(_04908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04944_));
 sky130_fd_sc_hd__o22a_1 _11085_ (.A1(\sha256cu.m_pad_pars.block_512[27][7] ),
    .A2(_04944_),
    .B1(_04753_),
    .B2(_04907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04945_));
 sky130_fd_sc_hd__o22a_1 _11086_ (.A1(_04753_),
    .A2(_04933_),
    .B1(_04788_),
    .B2(\sha256cu.m_pad_pars.block_512[11][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04946_));
 sky130_fd_sc_hd__inv_2 _11087_ (.A(_04784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04947_));
 sky130_fd_sc_hd__a32o_1 _11088_ (.A1(_04755_),
    .A2(_04756_),
    .A3(_04945_),
    .B1(_04946_),
    .B2(_04947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04948_));
 sky130_fd_sc_hd__a31o_1 _11089_ (.A1(_04756_),
    .A2(_04764_),
    .A3(_04943_),
    .B1(_04948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04949_));
 sky130_fd_sc_hd__a311o_1 _11090_ (.A1(_04736_),
    .A2(_04764_),
    .A3(_04932_),
    .B1(_04941_),
    .C1(_04949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04950_));
 sky130_fd_sc_hd__o221a_1 _11091_ (.A1(\sha256cu.data_in_padd[7] ),
    .A2(_04840_),
    .B1(_04931_),
    .B2(_04950_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00870_));
 sky130_fd_sc_hd__and2b_1 _11092_ (.A_N(\sha256cu.m_pad_pars.add_out2[3] ),
    .B(\sha256cu.m_pad_pars.add_out2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04951_));
 sky130_fd_sc_hd__or3b_1 _11093_ (.A(_04725_),
    .B(_04721_),
    .C_N(_04951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04952_));
 sky130_fd_sc_hd__or2b_1 _11094_ (.A(\sha256cu.m_pad_pars.add_512_block[1] ),
    .B_N(_01939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04953_));
 sky130_fd_sc_hd__or2_4 _11095_ (.A(_01953_),
    .B(_04953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04954_));
 sky130_fd_sc_hd__nor2_1 _11096_ (.A(_04771_),
    .B(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04955_));
 sky130_fd_sc_hd__o21bai_2 _11097_ (.A1(_04769_),
    .A2(_04954_),
    .B1_N(_04955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04956_));
 sky130_fd_sc_hd__nor2_4 _11098_ (.A(_04952_),
    .B(_04956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04957_));
 sky130_fd_sc_hd__and2b_1 _11099_ (.A_N(\sha256cu.m_pad_pars.add_out2[2] ),
    .B(\sha256cu.m_pad_pars.add_out2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04958_));
 sky130_fd_sc_hd__or3b_2 _11100_ (.A(_04725_),
    .B(_04721_),
    .C_N(_04958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04959_));
 sky130_fd_sc_hd__or2_4 _11101_ (.A(_04749_),
    .B(_04953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04960_));
 sky130_fd_sc_hd__o21a_1 _11102_ (.A1(_04701_),
    .A2(_04753_),
    .B1(_04960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04961_));
 sky130_fd_sc_hd__nor2_1 _11103_ (.A(_04769_),
    .B(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04962_));
 sky130_fd_sc_hd__nor2_4 _11104_ (.A(_04959_),
    .B(_04962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04963_));
 sky130_fd_sc_hd__o211a_2 _11105_ (.A1(_04907_),
    .A2(_04961_),
    .B1(_04958_),
    .C1(_04726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04964_));
 sky130_fd_sc_hd__a22o_1 _11106_ (.A1(\sha256cu.m_pad_pars.block_512[10][0] ),
    .A2(_04963_),
    .B1(_04964_),
    .B2(\sha256cu.m_pad_pars.block_512[26][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04965_));
 sky130_fd_sc_hd__or2b_1 _11107_ (.A(\sha256cu.m_pad_pars.add_out2[4] ),
    .B_N(\sha256cu.m_pad_pars.add_out2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04966_));
 sky130_fd_sc_hd__inv_2 _11108_ (.A(_04966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04967_));
 sky130_fd_sc_hd__nand2_1 _11109_ (.A(_04951_),
    .B(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04968_));
 sky130_fd_sc_hd__or2_2 _11110_ (.A(_04704_),
    .B(_04954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04969_));
 sky130_fd_sc_hd__inv_2 _11111_ (.A(_04797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04970_));
 sky130_fd_sc_hd__a2bb2o_2 _11112_ (.A1_N(_04791_),
    .A2_N(_04969_),
    .B1(_04970_),
    .B2(_04698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04971_));
 sky130_fd_sc_hd__nor2_4 _11113_ (.A(_04968_),
    .B(_04971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04972_));
 sky130_fd_sc_hd__nor2_2 _11114_ (.A(_04776_),
    .B(_04953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04973_));
 sky130_fd_sc_hd__nor2_1 _11115_ (.A(_04701_),
    .B(_04779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04974_));
 sky130_fd_sc_hd__nor2_2 _11116_ (.A(_04973_),
    .B(_04974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04975_));
 sky130_fd_sc_hd__nor2_1 _11117_ (.A(_04720_),
    .B(_04966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04976_));
 sky130_fd_sc_hd__o21a_2 _11118_ (.A1(_04913_),
    .A2(_04975_),
    .B1(_04976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04977_));
 sky130_fd_sc_hd__and3_1 _11119_ (.A(_04725_),
    .B(_04721_),
    .C(_04951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04978_));
 sky130_fd_sc_hd__or2_1 _11120_ (.A(_01952_),
    .B(_04969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04979_));
 sky130_fd_sc_hd__or2_1 _11121_ (.A(_04796_),
    .B(_04824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04980_));
 sky130_fd_sc_hd__and3_2 _11122_ (.A(_04978_),
    .B(_04979_),
    .C(_04980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04981_));
 sky130_fd_sc_hd__and3_2 _11123_ (.A(_04725_),
    .B(\sha256cu.m_pad_pars.add_out2[4] ),
    .C(_04958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04982_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(\sha256cu.m_pad_pars.m_size[8] ),
    .A1(\sha256cu.m_pad_pars.block_512[62][0] ),
    .S(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04983_));
 sky130_fd_sc_hd__and4_2 _11125_ (.A(\sha256cu.m_pad_pars.add_out2[5] ),
    .B(\sha256cu.m_pad_pars.add_out2[4] ),
    .C(\sha256cu.m_pad_pars.add_out2[3] ),
    .D(\sha256cu.m_pad_pars.add_out2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04984_));
 sky130_fd_sc_hd__a32o_1 _11126_ (.A1(\sha256cu.m_pad_pars.block_512[58][0] ),
    .A2(_01920_),
    .A3(_04982_),
    .B1(_04983_),
    .B2(_04984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04985_));
 sky130_fd_sc_hd__a221o_1 _11127_ (.A1(\sha256cu.m_pad_pars.block_512[46][0] ),
    .A2(_04977_),
    .B1(_04981_),
    .B2(\sha256cu.m_pad_pars.block_512[54][0] ),
    .C1(_04985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04986_));
 sky130_fd_sc_hd__or3_2 _11128_ (.A(_04725_),
    .B(_04721_),
    .C(_04720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04987_));
 sky130_fd_sc_hd__nor2_1 _11129_ (.A(_04769_),
    .B(_04975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04988_));
 sky130_fd_sc_hd__nor2_4 _11130_ (.A(_04987_),
    .B(_04988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04989_));
 sky130_fd_sc_hd__nor2_2 _11131_ (.A(\sha256cu.m_pad_pars.add_out2[3] ),
    .B(\sha256cu.m_pad_pars.add_out2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04990_));
 sky130_fd_sc_hd__nand2_2 _11132_ (.A(_04990_),
    .B(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04991_));
 sky130_fd_sc_hd__or2_1 _11133_ (.A(_01940_),
    .B(_04953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04992_));
 sky130_fd_sc_hd__buf_2 _11134_ (.A(_04992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04993_));
 sky130_fd_sc_hd__o21a_1 _11135_ (.A1(_04701_),
    .A2(_04758_),
    .B1(_04993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04994_));
 sky130_fd_sc_hd__nor2_1 _11136_ (.A(_04913_),
    .B(_04994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04995_));
 sky130_fd_sc_hd__nor2_4 _11137_ (.A(_04991_),
    .B(_04995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04996_));
 sky130_fd_sc_hd__or4_2 _11138_ (.A(_04725_),
    .B(_04721_),
    .C(\sha256cu.m_pad_pars.add_out2[3] ),
    .D(\sha256cu.m_pad_pars.add_out2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04997_));
 sky130_fd_sc_hd__nor2_1 _11139_ (.A(_04768_),
    .B(_04994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04998_));
 sky130_fd_sc_hd__nor2_2 _11140_ (.A(_04997_),
    .B(_04998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04999_));
 sky130_fd_sc_hd__or2_1 _11141_ (.A(_04912_),
    .B(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05000_));
 sky130_fd_sc_hd__and4b_4 _11142_ (.A_N(_04721_),
    .B(_04958_),
    .C(_05000_),
    .D(_04725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05001_));
 sky130_fd_sc_hd__a22o_1 _11143_ (.A1(\sha256cu.m_pad_pars.block_512[2][0] ),
    .A2(_04999_),
    .B1(_05001_),
    .B2(\sha256cu.m_pad_pars.block_512[42][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05002_));
 sky130_fd_sc_hd__a221o_1 _11144_ (.A1(\sha256cu.m_pad_pars.block_512[14][0] ),
    .A2(_04989_),
    .B1(_04996_),
    .B2(\sha256cu.m_pad_pars.block_512[34][0] ),
    .C1(_05002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05003_));
 sky130_fd_sc_hd__or2_2 _11145_ (.A(_04704_),
    .B(_04993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05004_));
 sky130_fd_sc_hd__nor2_1 _11146_ (.A(_04759_),
    .B(_04824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05005_));
 sky130_fd_sc_hd__o21bai_2 _11147_ (.A1(_01952_),
    .A2(_05004_),
    .B1_N(_05005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05006_));
 sky130_fd_sc_hd__inv_2 _11148_ (.A(_05006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05007_));
 sky130_fd_sc_hd__and4_4 _11149_ (.A(_04725_),
    .B(_04721_),
    .C(_04990_),
    .D(_05007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05008_));
 sky130_fd_sc_hd__o21a_2 _11150_ (.A1(_04747_),
    .A2(_04975_),
    .B1(_04727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05009_));
 sky130_fd_sc_hd__nand2_1 _11151_ (.A(_04699_),
    .B(_04925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05010_));
 sky130_fd_sc_hd__nor2_2 _11152_ (.A(_04771_),
    .B(_05010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05011_));
 sky130_fd_sc_hd__nor2_2 _11153_ (.A(_04746_),
    .B(_04954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05012_));
 sky130_fd_sc_hd__and4bb_2 _11154_ (.A_N(_05011_),
    .B_N(_05012_),
    .C(_04726_),
    .D(_04951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05013_));
 sky130_fd_sc_hd__o211a_2 _11155_ (.A1(_04747_),
    .A2(_04994_),
    .B1(_04990_),
    .C1(_04726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05014_));
 sky130_fd_sc_hd__a22o_1 _11156_ (.A1(\sha256cu.m_pad_pars.block_512[22][0] ),
    .A2(_05013_),
    .B1(_05014_),
    .B2(\sha256cu.m_pad_pars.block_512[18][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05015_));
 sky130_fd_sc_hd__a221o_1 _11157_ (.A1(\sha256cu.m_pad_pars.block_512[50][0] ),
    .A2(_05008_),
    .B1(_05009_),
    .B2(\sha256cu.m_pad_pars.block_512[30][0] ),
    .C1(_05015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05016_));
 sky130_fd_sc_hd__a2111o_1 _11158_ (.A1(\sha256cu.m_pad_pars.block_512[38][0] ),
    .A2(_04972_),
    .B1(_04986_),
    .C1(_05003_),
    .D1(_05016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05017_));
 sky130_fd_sc_hd__a211o_1 _11159_ (.A1(\sha256cu.m_pad_pars.block_512[6][0] ),
    .A2(_04957_),
    .B1(_04965_),
    .C1(_05017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05018_));
 sky130_fd_sc_hd__a22o_1 _11160_ (.A1(\sha256cu.data_in_padd[8] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00871_));
 sky130_fd_sc_hd__a22o_1 _11161_ (.A1(\sha256cu.m_pad_pars.block_512[6][1] ),
    .A2(_04957_),
    .B1(_04964_),
    .B2(\sha256cu.m_pad_pars.block_512[26][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05019_));
 sky130_fd_sc_hd__a22o_1 _11162_ (.A1(\sha256cu.m_pad_pars.block_512[2][1] ),
    .A2(_04999_),
    .B1(_04996_),
    .B2(\sha256cu.m_pad_pars.block_512[34][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05020_));
 sky130_fd_sc_hd__a221o_1 _11163_ (.A1(\sha256cu.m_pad_pars.block_512[10][1] ),
    .A2(_04963_),
    .B1(_04972_),
    .B2(\sha256cu.m_pad_pars.block_512[38][1] ),
    .C1(_05020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05021_));
 sky130_fd_sc_hd__a22o_1 _11164_ (.A1(\sha256cu.m_pad_pars.block_512[18][1] ),
    .A2(_05014_),
    .B1(_05009_),
    .B2(\sha256cu.m_pad_pars.block_512[30][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05022_));
 sky130_fd_sc_hd__a221o_1 _11165_ (.A1(\sha256cu.m_pad_pars.block_512[22][1] ),
    .A2(_05013_),
    .B1(_04977_),
    .B2(\sha256cu.m_pad_pars.block_512[46][1] ),
    .C1(_05022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05023_));
 sky130_fd_sc_hd__buf_4 _11166_ (.A(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05024_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(\sha256cu.m_pad_pars.m_size[9] ),
    .A1(\sha256cu.m_pad_pars.block_512[62][1] ),
    .S(_05024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05025_));
 sky130_fd_sc_hd__a32o_1 _11168_ (.A1(\sha256cu.m_pad_pars.block_512[58][1] ),
    .A2(_01921_),
    .A3(_04982_),
    .B1(_05025_),
    .B2(_04984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05026_));
 sky130_fd_sc_hd__a221o_1 _11169_ (.A1(\sha256cu.m_pad_pars.block_512[50][1] ),
    .A2(_05008_),
    .B1(_04981_),
    .B2(\sha256cu.m_pad_pars.block_512[54][1] ),
    .C1(_05026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05027_));
 sky130_fd_sc_hd__a2111o_1 _11170_ (.A1(\sha256cu.m_pad_pars.block_512[42][1] ),
    .A2(_05001_),
    .B1(_05021_),
    .C1(_05023_),
    .D1(_05027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05028_));
 sky130_fd_sc_hd__a211o_1 _11171_ (.A1(\sha256cu.m_pad_pars.block_512[14][1] ),
    .A2(_04989_),
    .B1(_05019_),
    .C1(_05028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05029_));
 sky130_fd_sc_hd__a22o_1 _11172_ (.A1(\sha256cu.data_in_padd[9] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00872_));
 sky130_fd_sc_hd__a22o_1 _11173_ (.A1(\sha256cu.m_pad_pars.block_512[62][2] ),
    .A2(_04984_),
    .B1(_04982_),
    .B2(\sha256cu.m_pad_pars.block_512[58][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05030_));
 sky130_fd_sc_hd__a22o_1 _11174_ (.A1(\sha256cu.m_pad_pars.block_512[2][2] ),
    .A2(_04999_),
    .B1(_05030_),
    .B2(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05031_));
 sky130_fd_sc_hd__a221o_1 _11175_ (.A1(\sha256cu.m_pad_pars.block_512[6][2] ),
    .A2(_04957_),
    .B1(_04989_),
    .B2(\sha256cu.m_pad_pars.block_512[14][2] ),
    .C1(_05031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05032_));
 sky130_fd_sc_hd__a22o_1 _11176_ (.A1(\sha256cu.m_pad_pars.block_512[26][2] ),
    .A2(_04964_),
    .B1(_05014_),
    .B2(\sha256cu.m_pad_pars.block_512[18][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05033_));
 sky130_fd_sc_hd__a221o_1 _11177_ (.A1(\sha256cu.m_pad_pars.block_512[10][2] ),
    .A2(_04963_),
    .B1(_05001_),
    .B2(\sha256cu.m_pad_pars.block_512[42][2] ),
    .C1(_05033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05034_));
 sky130_fd_sc_hd__a22o_1 _11178_ (.A1(\sha256cu.m_pad_pars.block_512[30][2] ),
    .A2(_05009_),
    .B1(_04977_),
    .B2(\sha256cu.m_pad_pars.block_512[46][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05035_));
 sky130_fd_sc_hd__or3_1 _11179_ (.A(_05032_),
    .B(_05034_),
    .C(_05035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05036_));
 sky130_fd_sc_hd__a22o_1 _11180_ (.A1(\sha256cu.m_pad_pars.block_512[34][2] ),
    .A2(_04996_),
    .B1(_04981_),
    .B2(\sha256cu.m_pad_pars.block_512[54][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05037_));
 sky130_fd_sc_hd__a221o_1 _11181_ (.A1(\sha256cu.m_pad_pars.block_512[50][2] ),
    .A2(_05008_),
    .B1(_04972_),
    .B2(\sha256cu.m_pad_pars.block_512[38][2] ),
    .C1(_05037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05038_));
 sky130_fd_sc_hd__a211o_1 _11182_ (.A1(\sha256cu.m_pad_pars.block_512[22][2] ),
    .A2(_05013_),
    .B1(_05038_),
    .C1(_01971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05039_));
 sky130_fd_sc_hd__buf_4 _11183_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05040_));
 sky130_fd_sc_hd__o221a_1 _11184_ (.A1(\sha256cu.data_in_padd[10] ),
    .A2(_04840_),
    .B1(_05036_),
    .B2(_05039_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00873_));
 sky130_fd_sc_hd__a22o_1 _11185_ (.A1(\sha256cu.m_pad_pars.block_512[30][3] ),
    .A2(_05009_),
    .B1(_04977_),
    .B2(\sha256cu.m_pad_pars.block_512[46][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05041_));
 sky130_fd_sc_hd__a22o_1 _11186_ (.A1(\sha256cu.m_pad_pars.block_512[62][3] ),
    .A2(_04984_),
    .B1(_04982_),
    .B2(\sha256cu.m_pad_pars.block_512[58][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05042_));
 sky130_fd_sc_hd__a22o_1 _11187_ (.A1(\sha256cu.m_pad_pars.block_512[2][3] ),
    .A2(_04999_),
    .B1(_05042_),
    .B2(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05043_));
 sky130_fd_sc_hd__a221o_1 _11188_ (.A1(\sha256cu.m_pad_pars.block_512[6][3] ),
    .A2(_04957_),
    .B1(_04989_),
    .B2(\sha256cu.m_pad_pars.block_512[14][3] ),
    .C1(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05044_));
 sky130_fd_sc_hd__a22o_1 _11189_ (.A1(\sha256cu.m_pad_pars.block_512[26][3] ),
    .A2(_04964_),
    .B1(_05014_),
    .B2(\sha256cu.m_pad_pars.block_512[18][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05045_));
 sky130_fd_sc_hd__a221o_1 _11190_ (.A1(\sha256cu.m_pad_pars.block_512[10][3] ),
    .A2(_04963_),
    .B1(_05001_),
    .B2(\sha256cu.m_pad_pars.block_512[42][3] ),
    .C1(_05045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05046_));
 sky130_fd_sc_hd__or3_1 _11191_ (.A(_05041_),
    .B(_05044_),
    .C(_05046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05047_));
 sky130_fd_sc_hd__a22o_1 _11192_ (.A1(\sha256cu.m_pad_pars.block_512[34][3] ),
    .A2(_04996_),
    .B1(_04981_),
    .B2(\sha256cu.m_pad_pars.block_512[54][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05048_));
 sky130_fd_sc_hd__a221o_1 _11193_ (.A1(\sha256cu.m_pad_pars.block_512[50][3] ),
    .A2(_05008_),
    .B1(_04972_),
    .B2(\sha256cu.m_pad_pars.block_512[38][3] ),
    .C1(_05048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05049_));
 sky130_fd_sc_hd__a211o_1 _11194_ (.A1(\sha256cu.m_pad_pars.block_512[22][3] ),
    .A2(_05013_),
    .B1(_05049_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05050_));
 sky130_fd_sc_hd__o221a_1 _11195_ (.A1(\sha256cu.data_in_padd[11] ),
    .A2(_04840_),
    .B1(_05047_),
    .B2(_05050_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00874_));
 sky130_fd_sc_hd__a22o_1 _11196_ (.A1(\sha256cu.m_pad_pars.block_512[26][4] ),
    .A2(_04964_),
    .B1(_05014_),
    .B2(\sha256cu.m_pad_pars.block_512[18][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05051_));
 sky130_fd_sc_hd__a22o_1 _11197_ (.A1(\sha256cu.m_pad_pars.block_512[62][4] ),
    .A2(_04984_),
    .B1(_04982_),
    .B2(\sha256cu.m_pad_pars.block_512[58][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05052_));
 sky130_fd_sc_hd__a22o_1 _11198_ (.A1(\sha256cu.m_pad_pars.block_512[2][4] ),
    .A2(_04999_),
    .B1(_05052_),
    .B2(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05053_));
 sky130_fd_sc_hd__a22o_1 _11199_ (.A1(\sha256cu.m_pad_pars.block_512[42][4] ),
    .A2(_05001_),
    .B1(_04989_),
    .B2(\sha256cu.m_pad_pars.block_512[14][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05054_));
 sky130_fd_sc_hd__a211o_1 _11200_ (.A1(\sha256cu.m_pad_pars.block_512[6][4] ),
    .A2(_04957_),
    .B1(_05053_),
    .C1(_05054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05055_));
 sky130_fd_sc_hd__a211o_1 _11201_ (.A1(\sha256cu.m_pad_pars.block_512[10][4] ),
    .A2(_04963_),
    .B1(_05051_),
    .C1(_05055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05056_));
 sky130_fd_sc_hd__a221o_1 _11202_ (.A1(\sha256cu.m_pad_pars.block_512[30][4] ),
    .A2(_05009_),
    .B1(_04977_),
    .B2(\sha256cu.m_pad_pars.block_512[46][4] ),
    .C1(_05056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05057_));
 sky130_fd_sc_hd__a22o_1 _11203_ (.A1(\sha256cu.m_pad_pars.block_512[34][4] ),
    .A2(_04996_),
    .B1(_04981_),
    .B2(\sha256cu.m_pad_pars.block_512[54][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05058_));
 sky130_fd_sc_hd__a221o_1 _11204_ (.A1(\sha256cu.m_pad_pars.block_512[50][4] ),
    .A2(_05008_),
    .B1(_04972_),
    .B2(\sha256cu.m_pad_pars.block_512[38][4] ),
    .C1(_05058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05059_));
 sky130_fd_sc_hd__a211o_1 _11205_ (.A1(\sha256cu.m_pad_pars.block_512[22][4] ),
    .A2(_05013_),
    .B1(_05059_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05060_));
 sky130_fd_sc_hd__o221a_1 _11206_ (.A1(\sha256cu.data_in_padd[12] ),
    .A2(_04840_),
    .B1(_05057_),
    .B2(_05060_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00875_));
 sky130_fd_sc_hd__a22o_1 _11207_ (.A1(\sha256cu.m_pad_pars.block_512[26][5] ),
    .A2(_04964_),
    .B1(_05014_),
    .B2(\sha256cu.m_pad_pars.block_512[18][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05061_));
 sky130_fd_sc_hd__a22o_1 _11208_ (.A1(\sha256cu.m_pad_pars.block_512[62][5] ),
    .A2(_04984_),
    .B1(_04982_),
    .B2(\sha256cu.m_pad_pars.block_512[58][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05062_));
 sky130_fd_sc_hd__and2_1 _11209_ (.A(_05024_),
    .B(_05062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05063_));
 sky130_fd_sc_hd__a221o_1 _11210_ (.A1(\sha256cu.m_pad_pars.block_512[2][5] ),
    .A2(_04999_),
    .B1(_04989_),
    .B2(\sha256cu.m_pad_pars.block_512[14][5] ),
    .C1(_05063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05064_));
 sky130_fd_sc_hd__a221o_1 _11211_ (.A1(\sha256cu.m_pad_pars.block_512[6][5] ),
    .A2(_04957_),
    .B1(_05001_),
    .B2(\sha256cu.m_pad_pars.block_512[42][5] ),
    .C1(_05064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05065_));
 sky130_fd_sc_hd__a211o_1 _11212_ (.A1(\sha256cu.m_pad_pars.block_512[10][5] ),
    .A2(_04963_),
    .B1(_05061_),
    .C1(_05065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05066_));
 sky130_fd_sc_hd__a221o_1 _11213_ (.A1(\sha256cu.m_pad_pars.block_512[30][5] ),
    .A2(_05009_),
    .B1(_04977_),
    .B2(\sha256cu.m_pad_pars.block_512[46][5] ),
    .C1(_05066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05067_));
 sky130_fd_sc_hd__a22o_1 _11214_ (.A1(\sha256cu.m_pad_pars.block_512[34][5] ),
    .A2(_04996_),
    .B1(_04981_),
    .B2(\sha256cu.m_pad_pars.block_512[54][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05068_));
 sky130_fd_sc_hd__a221o_1 _11215_ (.A1(\sha256cu.m_pad_pars.block_512[50][5] ),
    .A2(_05008_),
    .B1(_04972_),
    .B2(\sha256cu.m_pad_pars.block_512[38][5] ),
    .C1(_05068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05069_));
 sky130_fd_sc_hd__a211o_1 _11216_ (.A1(\sha256cu.m_pad_pars.block_512[22][5] ),
    .A2(_05013_),
    .B1(_05069_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05070_));
 sky130_fd_sc_hd__o221a_1 _11217_ (.A1(\sha256cu.data_in_padd[13] ),
    .A2(_04840_),
    .B1(_05067_),
    .B2(_05070_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00876_));
 sky130_fd_sc_hd__a22o_1 _11218_ (.A1(\sha256cu.m_pad_pars.block_512[2][6] ),
    .A2(_04999_),
    .B1(_04972_),
    .B2(\sha256cu.m_pad_pars.block_512[38][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05071_));
 sky130_fd_sc_hd__a221o_1 _11219_ (.A1(\sha256cu.m_pad_pars.block_512[6][6] ),
    .A2(_04957_),
    .B1(_04989_),
    .B2(\sha256cu.m_pad_pars.block_512[14][6] ),
    .C1(_05071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05072_));
 sky130_fd_sc_hd__a22o_1 _11220_ (.A1(\sha256cu.m_pad_pars.block_512[62][6] ),
    .A2(_04984_),
    .B1(_04982_),
    .B2(\sha256cu.m_pad_pars.block_512[58][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05073_));
 sky130_fd_sc_hd__and2_1 _11221_ (.A(_05024_),
    .B(_05073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05074_));
 sky130_fd_sc_hd__a221o_1 _11222_ (.A1(\sha256cu.m_pad_pars.block_512[46][6] ),
    .A2(_04977_),
    .B1(_04981_),
    .B2(\sha256cu.m_pad_pars.block_512[54][6] ),
    .C1(_05074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05075_));
 sky130_fd_sc_hd__a221o_1 _11223_ (.A1(\sha256cu.m_pad_pars.block_512[26][6] ),
    .A2(_04964_),
    .B1(_05009_),
    .B2(\sha256cu.m_pad_pars.block_512[30][6] ),
    .C1(_05075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05076_));
 sky130_fd_sc_hd__a211o_1 _11224_ (.A1(\sha256cu.m_pad_pars.block_512[50][6] ),
    .A2(_05008_),
    .B1(_05072_),
    .C1(_05076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05077_));
 sky130_fd_sc_hd__a221o_1 _11225_ (.A1(\sha256cu.m_pad_pars.block_512[10][6] ),
    .A2(_04963_),
    .B1(_04996_),
    .B2(\sha256cu.m_pad_pars.block_512[34][6] ),
    .C1(_05077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05078_));
 sky130_fd_sc_hd__a22o_1 _11226_ (.A1(\sha256cu.m_pad_pars.block_512[42][6] ),
    .A2(_05001_),
    .B1(_05013_),
    .B2(\sha256cu.m_pad_pars.block_512[22][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05079_));
 sky130_fd_sc_hd__a211o_1 _11227_ (.A1(\sha256cu.m_pad_pars.block_512[18][6] ),
    .A2(_05014_),
    .B1(_05079_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05080_));
 sky130_fd_sc_hd__o221a_1 _11228_ (.A1(\sha256cu.data_in_padd[14] ),
    .A2(_04840_),
    .B1(_05078_),
    .B2(_05080_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00877_));
 sky130_fd_sc_hd__buf_4 _11229_ (.A(_04907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05081_));
 sky130_fd_sc_hd__a31o_1 _11230_ (.A1(_04698_),
    .A2(_04908_),
    .A3(_04785_),
    .B1(\sha256cu.m_pad_pars.block_512[26][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05082_));
 sky130_fd_sc_hd__o21a_1 _11231_ (.A1(_05081_),
    .A2(_04960_),
    .B1(_05082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05083_));
 sky130_fd_sc_hd__a21o_1 _11232_ (.A1(_04698_),
    .A2(_04970_),
    .B1(\sha256cu.m_pad_pars.block_512[38][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05084_));
 sky130_fd_sc_hd__o21a_1 _11233_ (.A1(_04917_),
    .A2(_04954_),
    .B1(_05084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05085_));
 sky130_fd_sc_hd__nor2_1 _11234_ (.A(_04753_),
    .B(_04794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05086_));
 sky130_fd_sc_hd__o22a_1 _11235_ (.A1(_04913_),
    .A2(_04960_),
    .B1(_05086_),
    .B2(\sha256cu.m_pad_pars.block_512[42][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05087_));
 sky130_fd_sc_hd__and3_1 _11236_ (.A(_04958_),
    .B(_04967_),
    .C(_05087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05088_));
 sky130_fd_sc_hd__a31o_1 _11237_ (.A1(_04951_),
    .A2(_04967_),
    .A3(_05085_),
    .B1(_05088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05089_));
 sky130_fd_sc_hd__and3_1 _11238_ (.A(_04698_),
    .B(_04785_),
    .C(_04786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05090_));
 sky130_fd_sc_hd__or2_1 _11239_ (.A(_04768_),
    .B(_04960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05091_));
 sky130_fd_sc_hd__inv_2 _11240_ (.A(_04959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05092_));
 sky130_fd_sc_hd__o211a_1 _11241_ (.A1(\sha256cu.m_pad_pars.block_512[10][7] ),
    .A2(_05090_),
    .B1(_05091_),
    .C1(_05092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05093_));
 sky130_fd_sc_hd__a311o_1 _11242_ (.A1(_04726_),
    .A2(_04958_),
    .A3(_05083_),
    .B1(_05089_),
    .C1(_05093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_1 _11243_ (.A(_04702_),
    .B(_04780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _11244_ (.A(_04786_),
    .B(_04973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05096_));
 sky130_fd_sc_hd__o21a_1 _11245_ (.A1(\sha256cu.m_pad_pars.block_512[14][7] ),
    .A2(_05095_),
    .B1(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05097_));
 sky130_fd_sc_hd__and2b_1 _11246_ (.A_N(_04987_),
    .B(_05097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05098_));
 sky130_fd_sc_hd__o22a_1 _11247_ (.A1(\sha256cu.m_pad_pars.block_512[6][7] ),
    .A2(_04955_),
    .B1(_04954_),
    .B2(_04933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05099_));
 sky130_fd_sc_hd__and2b_1 _11248_ (.A_N(_04952_),
    .B(_05099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05100_));
 sky130_fd_sc_hd__nand2_1 _11249_ (.A(_04908_),
    .B(_04973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05101_));
 sky130_fd_sc_hd__a22o_1 _11250_ (.A1(_04908_),
    .A2(_04974_),
    .B1(_05101_),
    .B2(\sha256cu.m_pad_pars.block_512[30][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05102_));
 sky130_fd_sc_hd__nor2_1 _11251_ (.A(_04796_),
    .B(_04824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05103_));
 sky130_fd_sc_hd__o21a_1 _11252_ (.A1(\sha256cu.m_pad_pars.block_512[54][7] ),
    .A2(_05103_),
    .B1(_04979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05104_));
 sky130_fd_sc_hd__a22o_1 _11253_ (.A1(\sha256cu.m_pad_pars.block_512[62][7] ),
    .A2(_04984_),
    .B1(_04982_),
    .B2(\sha256cu.m_pad_pars.block_512[58][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05105_));
 sky130_fd_sc_hd__a22o_1 _11254_ (.A1(_04978_),
    .A2(_05104_),
    .B1(_05105_),
    .B2(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05106_));
 sky130_fd_sc_hd__nor2_1 _11255_ (.A(_04759_),
    .B(_04807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05107_));
 sky130_fd_sc_hd__o22a_1 _11256_ (.A1(_04747_),
    .A2(_04993_),
    .B1(_05107_),
    .B2(\sha256cu.m_pad_pars.block_512[18][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05108_));
 sky130_fd_sc_hd__o22a_1 _11257_ (.A1(_01952_),
    .A2(_05004_),
    .B1(_05005_),
    .B2(\sha256cu.m_pad_pars.block_512[50][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05109_));
 sky130_fd_sc_hd__and4_1 _11258_ (.A(_04725_),
    .B(_04721_),
    .C(_04990_),
    .D(_05109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05110_));
 sky130_fd_sc_hd__o21ba_1 _11259_ (.A1(\sha256cu.m_pad_pars.block_512[22][7] ),
    .A2(_05011_),
    .B1_N(_05012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05111_));
 sky130_fd_sc_hd__nand2_1 _11260_ (.A(_04801_),
    .B(_04973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05112_));
 sky130_fd_sc_hd__a22o_1 _11261_ (.A1(_04801_),
    .A2(_04974_),
    .B1(_05112_),
    .B2(\sha256cu.m_pad_pars.block_512[46][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05113_));
 sky130_fd_sc_hd__a32o_1 _11262_ (.A1(_04726_),
    .A2(_04951_),
    .A3(_05111_),
    .B1(_05113_),
    .B2(_04976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05114_));
 sky130_fd_sc_hd__a311o_1 _11263_ (.A1(_04726_),
    .A2(_04990_),
    .A3(_05108_),
    .B1(_05110_),
    .C1(_05114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05115_));
 sky130_fd_sc_hd__a2111o_1 _11264_ (.A1(_04727_),
    .A2(_05102_),
    .B1(_05106_),
    .C1(_05115_),
    .D1(_01969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05116_));
 sky130_fd_sc_hd__nor2_1 _11265_ (.A(_04702_),
    .B(_04758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05117_));
 sky130_fd_sc_hd__a31o_1 _11266_ (.A1(_01944_),
    .A2(_04699_),
    .A3(_05117_),
    .B1(\sha256cu.m_pad_pars.block_512[2][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05118_));
 sky130_fd_sc_hd__o21ai_1 _11267_ (.A1(_04933_),
    .A2(_04993_),
    .B1(_05118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05119_));
 sky130_fd_sc_hd__a21o_1 _11268_ (.A1(_04801_),
    .A2(_05117_),
    .B1(\sha256cu.m_pad_pars.block_512[34][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05120_));
 sky130_fd_sc_hd__o21ai_1 _11269_ (.A1(_04917_),
    .A2(_04993_),
    .B1(_05120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05121_));
 sky130_fd_sc_hd__o22a_1 _11270_ (.A1(_04997_),
    .A2(_05119_),
    .B1(_05121_),
    .B2(_04991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05122_));
 sky130_fd_sc_hd__or4b_1 _11271_ (.A(_05098_),
    .B(_05100_),
    .C(_05116_),
    .D_N(_05122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05123_));
 sky130_fd_sc_hd__o221a_1 _11272_ (.A1(\sha256cu.data_in_padd[15] ),
    .A2(_01963_),
    .B1(_05094_),
    .B2(_05123_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00878_));
 sky130_fd_sc_hd__a211o_2 _11273_ (.A1(_04702_),
    .A2(_01939_),
    .B1(_04776_),
    .C1(\sha256cu.m_pad_pars.add_512_block[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05124_));
 sky130_fd_sc_hd__nor2b_2 _11274_ (.A(\sha256cu.m_pad_pars.add_out1[4] ),
    .B_N(\sha256cu.m_pad_pars.add_out1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05125_));
 sky130_fd_sc_hd__o211a_2 _11275_ (.A1(_04913_),
    .A2(_05124_),
    .B1(_05125_),
    .C1(_01977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05126_));
 sky130_fd_sc_hd__nor2_2 _11276_ (.A(\sha256cu.m_pad_pars.add_out1[5] ),
    .B(\sha256cu.m_pad_pars.add_out1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05127_));
 sky130_fd_sc_hd__o211a_2 _11277_ (.A1(_04933_),
    .A2(_05124_),
    .B1(_05127_),
    .C1(_01977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05128_));
 sky130_fd_sc_hd__or2_2 _11278_ (.A(_01941_),
    .B(_04749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05129_));
 sky130_fd_sc_hd__o21a_1 _11279_ (.A1(_04702_),
    .A2(_04960_),
    .B1(_05129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05130_));
 sky130_fd_sc_hd__or2_1 _11280_ (.A(_04913_),
    .B(_05130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05131_));
 sky130_fd_sc_hd__and4b_2 _11281_ (.A_N(\sha256cu.m_pad_pars.add_out1[2] ),
    .B(_05125_),
    .C(_05131_),
    .D(\sha256cu.m_pad_pars.add_out1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05132_));
 sky130_fd_sc_hd__a22o_1 _11282_ (.A1(\sha256cu.m_pad_pars.block_512[13][0] ),
    .A2(_05128_),
    .B1(_05132_),
    .B2(\sha256cu.m_pad_pars.block_512[41][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05133_));
 sky130_fd_sc_hd__nor2_2 _11283_ (.A(\sha256cu.m_pad_pars.add_out1[3] ),
    .B(\sha256cu.m_pad_pars.add_out1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05134_));
 sky130_fd_sc_hd__o211a_2 _11284_ (.A1(_04787_),
    .A2(_04993_),
    .B1(_05127_),
    .C1(_05134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05135_));
 sky130_fd_sc_hd__nand2_4 _11285_ (.A(_01942_),
    .B(_04699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05136_));
 sky130_fd_sc_hd__o22a_1 _11286_ (.A1(_04807_),
    .A2(_05004_),
    .B1(_05136_),
    .B2(_04805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05137_));
 sky130_fd_sc_hd__and3_2 _11287_ (.A(_01985_),
    .B(_05134_),
    .C(_05137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05138_));
 sky130_fd_sc_hd__and2b_2 _11288_ (.A_N(\sha256cu.m_pad_pars.add_out1[2] ),
    .B(\sha256cu.m_pad_pars.add_out1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05139_));
 sky130_fd_sc_hd__o211a_2 _11289_ (.A1(_04747_),
    .A2(_05130_),
    .B1(_05139_),
    .C1(_01985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05140_));
 sky130_fd_sc_hd__o211a_2 _11290_ (.A1(_04747_),
    .A2(_05124_),
    .B1(_01977_),
    .C1(_01985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05141_));
 sky130_fd_sc_hd__a22o_1 _11291_ (.A1(\sha256cu.m_pad_pars.block_512[25][0] ),
    .A2(_05140_),
    .B1(_05141_),
    .B2(\sha256cu.m_pad_pars.block_512[29][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05142_));
 sky130_fd_sc_hd__a221o_1 _11292_ (.A1(\sha256cu.m_pad_pars.block_512[1][0] ),
    .A2(_05135_),
    .B1(_05138_),
    .B2(\sha256cu.m_pad_pars.block_512[17][0] ),
    .C1(_05142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05143_));
 sky130_fd_sc_hd__o211a_2 _11293_ (.A1(_04769_),
    .A2(_05130_),
    .B1(_05139_),
    .C1(_05127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05144_));
 sky130_fd_sc_hd__nor3_1 _11294_ (.A(_04705_),
    .B(_04792_),
    .C(_04993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05145_));
 sky130_fd_sc_hd__o21ba_1 _11295_ (.A1(_04819_),
    .A2(_05136_),
    .B1_N(_05145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05146_));
 sky130_fd_sc_hd__and3_2 _11296_ (.A(_05125_),
    .B(_05134_),
    .C(_05146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05147_));
 sky130_fd_sc_hd__a22o_1 _11297_ (.A1(\sha256cu.m_pad_pars.block_512[9][0] ),
    .A2(_05144_),
    .B1(_05147_),
    .B2(\sha256cu.m_pad_pars.block_512[33][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05148_));
 sky130_fd_sc_hd__and2_1 _11298_ (.A(\sha256cu.m_pad_pars.add_out1[5] ),
    .B(\sha256cu.m_pad_pars.add_out1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05149_));
 sky130_fd_sc_hd__and2_1 _11299_ (.A(_05134_),
    .B(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05150_));
 sky130_fd_sc_hd__o221a_2 _11300_ (.A1(_04824_),
    .A2(_05004_),
    .B1(_05136_),
    .B2(_01952_),
    .C1(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05151_));
 sky130_fd_sc_hd__nor2b_2 _11301_ (.A(\sha256cu.m_pad_pars.add_out1[3] ),
    .B_N(\sha256cu.m_pad_pars.add_out1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05152_));
 sky130_fd_sc_hd__or2_1 _11302_ (.A(_01941_),
    .B(_01953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05153_));
 sky130_fd_sc_hd__clkbuf_4 _11303_ (.A(_05153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05154_));
 sky130_fd_sc_hd__nor2_1 _11304_ (.A(_04807_),
    .B(_04969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05155_));
 sky130_fd_sc_hd__o21bai_1 _11305_ (.A1(_04746_),
    .A2(_05154_),
    .B1_N(_05155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05156_));
 sky130_fd_sc_hd__inv_1 _11306_ (.A(_05156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05157_));
 sky130_fd_sc_hd__and3_2 _11307_ (.A(_01985_),
    .B(_05152_),
    .C(_05157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05158_));
 sky130_fd_sc_hd__o22a_2 _11308_ (.A1(\sha256cu.m_pad_pars.temp_chk ),
    .A2(_04954_),
    .B1(_05154_),
    .B2(\sha256cu.m_pad_pars.add_512_block[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05159_));
 sky130_fd_sc_hd__o211a_2 _11309_ (.A1(_04768_),
    .A2(_05159_),
    .B1(_05152_),
    .C1(_05127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05160_));
 sky130_fd_sc_hd__o311a_2 _11310_ (.A1(_01950_),
    .A2(_04704_),
    .A3(_05159_),
    .B1(_05149_),
    .C1(_05152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05161_));
 sky130_fd_sc_hd__and2_2 _11311_ (.A(_01977_),
    .B(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05162_));
 sky130_fd_sc_hd__and2_2 _11312_ (.A(_05139_),
    .B(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05163_));
 sky130_fd_sc_hd__a22o_1 _11313_ (.A1(\sha256cu.m_pad_pars.block_512[61][0] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05164_));
 sky130_fd_sc_hd__o211a_2 _11314_ (.A1(_04912_),
    .A2(_05159_),
    .B1(_05152_),
    .C1(_05125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05165_));
 sky130_fd_sc_hd__a22o_1 _11315_ (.A1(_05024_),
    .A2(_05164_),
    .B1(_05165_),
    .B2(\sha256cu.m_pad_pars.block_512[37][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05166_));
 sky130_fd_sc_hd__a221o_1 _11316_ (.A1(\sha256cu.m_pad_pars.block_512[5][0] ),
    .A2(_05160_),
    .B1(_05161_),
    .B2(\sha256cu.m_pad_pars.block_512[53][0] ),
    .C1(_05166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05167_));
 sky130_fd_sc_hd__a221o_1 _11317_ (.A1(\sha256cu.m_pad_pars.block_512[49][0] ),
    .A2(_05151_),
    .B1(_05158_),
    .B2(\sha256cu.m_pad_pars.block_512[21][0] ),
    .C1(_05167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05168_));
 sky130_fd_sc_hd__or3_1 _11318_ (.A(_05143_),
    .B(_05148_),
    .C(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05169_));
 sky130_fd_sc_hd__a211o_1 _11319_ (.A1(\sha256cu.m_pad_pars.block_512[45][0] ),
    .A2(_05126_),
    .B1(_05133_),
    .C1(_05169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05170_));
 sky130_fd_sc_hd__a22o_1 _11320_ (.A1(\sha256cu.data_in_padd[16] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00879_));
 sky130_fd_sc_hd__and2_1 _11321_ (.A(\sha256cu.m_pad_pars.block_512[45][1] ),
    .B(_05126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05171_));
 sky130_fd_sc_hd__a221o_1 _11322_ (.A1(\sha256cu.m_pad_pars.block_512[13][1] ),
    .A2(_05128_),
    .B1(_05132_),
    .B2(\sha256cu.m_pad_pars.block_512[41][1] ),
    .C1(_05171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05172_));
 sky130_fd_sc_hd__a22o_1 _11323_ (.A1(\sha256cu.m_pad_pars.block_512[1][1] ),
    .A2(_05135_),
    .B1(_05151_),
    .B2(\sha256cu.m_pad_pars.block_512[49][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05173_));
 sky130_fd_sc_hd__a221o_1 _11324_ (.A1(\sha256cu.m_pad_pars.block_512[29][1] ),
    .A2(_05141_),
    .B1(_05138_),
    .B2(\sha256cu.m_pad_pars.block_512[17][1] ),
    .C1(_05173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05174_));
 sky130_fd_sc_hd__a22o_1 _11325_ (.A1(\sha256cu.m_pad_pars.block_512[61][1] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05175_));
 sky130_fd_sc_hd__a22o_1 _11326_ (.A1(\sha256cu.m_pad_pars.block_512[53][1] ),
    .A2(_05161_),
    .B1(_05175_),
    .B2(_05024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05176_));
 sky130_fd_sc_hd__a221o_1 _11327_ (.A1(\sha256cu.m_pad_pars.block_512[5][1] ),
    .A2(_05160_),
    .B1(_05165_),
    .B2(\sha256cu.m_pad_pars.block_512[37][1] ),
    .C1(_05176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05177_));
 sky130_fd_sc_hd__a221o_1 _11328_ (.A1(\sha256cu.m_pad_pars.block_512[25][1] ),
    .A2(_05140_),
    .B1(_05158_),
    .B2(\sha256cu.m_pad_pars.block_512[21][1] ),
    .C1(_05177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05178_));
 sky130_fd_sc_hd__a221o_1 _11329_ (.A1(\sha256cu.m_pad_pars.block_512[9][1] ),
    .A2(_05144_),
    .B1(_05147_),
    .B2(\sha256cu.m_pad_pars.block_512[33][1] ),
    .C1(_05178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05179_));
 sky130_fd_sc_hd__or3_1 _11330_ (.A(_05172_),
    .B(_05174_),
    .C(_05179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05180_));
 sky130_fd_sc_hd__a22o_1 _11331_ (.A1(\sha256cu.data_in_padd[17] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00880_));
 sky130_fd_sc_hd__and2_1 _11332_ (.A(\sha256cu.m_pad_pars.block_512[45][2] ),
    .B(_05126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05181_));
 sky130_fd_sc_hd__a221o_1 _11333_ (.A1(\sha256cu.m_pad_pars.block_512[13][2] ),
    .A2(_05128_),
    .B1(_05132_),
    .B2(\sha256cu.m_pad_pars.block_512[41][2] ),
    .C1(_05181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05182_));
 sky130_fd_sc_hd__a22o_1 _11334_ (.A1(\sha256cu.m_pad_pars.block_512[1][2] ),
    .A2(_05135_),
    .B1(_05151_),
    .B2(\sha256cu.m_pad_pars.block_512[49][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05183_));
 sky130_fd_sc_hd__a221o_1 _11335_ (.A1(\sha256cu.m_pad_pars.block_512[17][2] ),
    .A2(_05138_),
    .B1(_05158_),
    .B2(\sha256cu.m_pad_pars.block_512[21][2] ),
    .C1(_05183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05184_));
 sky130_fd_sc_hd__a22o_1 _11336_ (.A1(\sha256cu.m_pad_pars.block_512[61][2] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05185_));
 sky130_fd_sc_hd__a22o_1 _11337_ (.A1(\sha256cu.m_pad_pars.block_512[37][2] ),
    .A2(_05165_),
    .B1(_05185_),
    .B2(_05024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05186_));
 sky130_fd_sc_hd__a221o_1 _11338_ (.A1(\sha256cu.m_pad_pars.block_512[5][2] ),
    .A2(_05160_),
    .B1(_05161_),
    .B2(\sha256cu.m_pad_pars.block_512[53][2] ),
    .C1(_05186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05187_));
 sky130_fd_sc_hd__a221o_1 _11339_ (.A1(\sha256cu.m_pad_pars.block_512[25][2] ),
    .A2(_05140_),
    .B1(_05141_),
    .B2(\sha256cu.m_pad_pars.block_512[29][2] ),
    .C1(_05187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05188_));
 sky130_fd_sc_hd__a221o_1 _11340_ (.A1(\sha256cu.m_pad_pars.block_512[9][2] ),
    .A2(_05144_),
    .B1(_05147_),
    .B2(\sha256cu.m_pad_pars.block_512[33][2] ),
    .C1(_05188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05189_));
 sky130_fd_sc_hd__or3_1 _11341_ (.A(_05182_),
    .B(_05184_),
    .C(_05189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05190_));
 sky130_fd_sc_hd__a22o_1 _11342_ (.A1(\sha256cu.data_in_padd[18] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00881_));
 sky130_fd_sc_hd__a22o_1 _11343_ (.A1(\sha256cu.m_pad_pars.block_512[13][3] ),
    .A2(_05128_),
    .B1(_05144_),
    .B2(\sha256cu.m_pad_pars.block_512[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05191_));
 sky130_fd_sc_hd__a21o_1 _11344_ (.A1(\sha256cu.m_pad_pars.block_512[33][3] ),
    .A2(_05147_),
    .B1(_05191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05192_));
 sky130_fd_sc_hd__a22o_1 _11345_ (.A1(\sha256cu.m_pad_pars.block_512[25][3] ),
    .A2(_05140_),
    .B1(_05138_),
    .B2(\sha256cu.m_pad_pars.block_512[17][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05193_));
 sky130_fd_sc_hd__a221o_1 _11346_ (.A1(\sha256cu.m_pad_pars.block_512[29][3] ),
    .A2(_05141_),
    .B1(_05135_),
    .B2(\sha256cu.m_pad_pars.block_512[1][3] ),
    .C1(_05193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05194_));
 sky130_fd_sc_hd__a22o_1 _11347_ (.A1(\sha256cu.m_pad_pars.block_512[61][3] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05195_));
 sky130_fd_sc_hd__a22o_1 _11348_ (.A1(\sha256cu.m_pad_pars.block_512[5][3] ),
    .A2(_05160_),
    .B1(_05195_),
    .B2(_05024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05196_));
 sky130_fd_sc_hd__a221o_1 _11349_ (.A1(\sha256cu.m_pad_pars.block_512[53][3] ),
    .A2(_05161_),
    .B1(_05165_),
    .B2(\sha256cu.m_pad_pars.block_512[37][3] ),
    .C1(_05196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05197_));
 sky130_fd_sc_hd__a221o_1 _11350_ (.A1(\sha256cu.m_pad_pars.block_512[49][3] ),
    .A2(_05151_),
    .B1(_05158_),
    .B2(\sha256cu.m_pad_pars.block_512[21][3] ),
    .C1(_05197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05198_));
 sky130_fd_sc_hd__a221o_1 _11351_ (.A1(\sha256cu.m_pad_pars.block_512[45][3] ),
    .A2(_05126_),
    .B1(_05132_),
    .B2(\sha256cu.m_pad_pars.block_512[41][3] ),
    .C1(_05198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05199_));
 sky130_fd_sc_hd__or3_1 _11352_ (.A(_05192_),
    .B(_05194_),
    .C(_05199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05200_));
 sky130_fd_sc_hd__a22o_1 _11353_ (.A1(\sha256cu.data_in_padd[19] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00882_));
 sky130_fd_sc_hd__and2_1 _11354_ (.A(\sha256cu.m_pad_pars.block_512[45][4] ),
    .B(_05126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05201_));
 sky130_fd_sc_hd__a221o_1 _11355_ (.A1(\sha256cu.m_pad_pars.block_512[13][4] ),
    .A2(_05128_),
    .B1(_05147_),
    .B2(\sha256cu.m_pad_pars.block_512[33][4] ),
    .C1(_05201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05202_));
 sky130_fd_sc_hd__a22o_1 _11356_ (.A1(\sha256cu.m_pad_pars.block_512[17][4] ),
    .A2(_05138_),
    .B1(_05151_),
    .B2(\sha256cu.m_pad_pars.block_512[49][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05203_));
 sky130_fd_sc_hd__a221o_1 _11357_ (.A1(\sha256cu.m_pad_pars.block_512[1][4] ),
    .A2(_05135_),
    .B1(_05158_),
    .B2(\sha256cu.m_pad_pars.block_512[21][4] ),
    .C1(_05203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05204_));
 sky130_fd_sc_hd__a22o_1 _11358_ (.A1(\sha256cu.m_pad_pars.block_512[61][4] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05205_));
 sky130_fd_sc_hd__a22o_1 _11359_ (.A1(\sha256cu.m_pad_pars.block_512[37][4] ),
    .A2(_05165_),
    .B1(_05205_),
    .B2(_05024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05206_));
 sky130_fd_sc_hd__a221o_1 _11360_ (.A1(\sha256cu.m_pad_pars.block_512[5][4] ),
    .A2(_05160_),
    .B1(_05161_),
    .B2(\sha256cu.m_pad_pars.block_512[53][4] ),
    .C1(_05206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05207_));
 sky130_fd_sc_hd__a221o_1 _11361_ (.A1(\sha256cu.m_pad_pars.block_512[25][4] ),
    .A2(_05140_),
    .B1(_05141_),
    .B2(\sha256cu.m_pad_pars.block_512[29][4] ),
    .C1(_05207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05208_));
 sky130_fd_sc_hd__a221o_1 _11362_ (.A1(\sha256cu.m_pad_pars.block_512[41][4] ),
    .A2(_05132_),
    .B1(_05144_),
    .B2(\sha256cu.m_pad_pars.block_512[9][4] ),
    .C1(_05208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05209_));
 sky130_fd_sc_hd__or3_1 _11363_ (.A(_05202_),
    .B(_05204_),
    .C(_05209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05210_));
 sky130_fd_sc_hd__a22o_1 _11364_ (.A1(\sha256cu.data_in_padd[20] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00883_));
 sky130_fd_sc_hd__and2_1 _11365_ (.A(\sha256cu.m_pad_pars.block_512[45][5] ),
    .B(_05126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05211_));
 sky130_fd_sc_hd__a221o_1 _11366_ (.A1(\sha256cu.m_pad_pars.block_512[13][5] ),
    .A2(_05128_),
    .B1(_05132_),
    .B2(\sha256cu.m_pad_pars.block_512[41][5] ),
    .C1(_05211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05212_));
 sky130_fd_sc_hd__a22o_1 _11367_ (.A1(\sha256cu.m_pad_pars.block_512[25][5] ),
    .A2(_05140_),
    .B1(_05141_),
    .B2(\sha256cu.m_pad_pars.block_512[29][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05213_));
 sky130_fd_sc_hd__a221o_1 _11368_ (.A1(\sha256cu.m_pad_pars.block_512[1][5] ),
    .A2(_05135_),
    .B1(_05138_),
    .B2(\sha256cu.m_pad_pars.block_512[17][5] ),
    .C1(_05213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05214_));
 sky130_fd_sc_hd__a22o_1 _11369_ (.A1(\sha256cu.m_pad_pars.block_512[61][5] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05215_));
 sky130_fd_sc_hd__a22o_1 _11370_ (.A1(\sha256cu.m_pad_pars.block_512[37][5] ),
    .A2(_05165_),
    .B1(_05215_),
    .B2(_05024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05216_));
 sky130_fd_sc_hd__a221o_1 _11371_ (.A1(\sha256cu.m_pad_pars.block_512[5][5] ),
    .A2(_05160_),
    .B1(_05161_),
    .B2(\sha256cu.m_pad_pars.block_512[53][5] ),
    .C1(_05216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05217_));
 sky130_fd_sc_hd__a221o_1 _11372_ (.A1(\sha256cu.m_pad_pars.block_512[49][5] ),
    .A2(_05151_),
    .B1(_05158_),
    .B2(\sha256cu.m_pad_pars.block_512[21][5] ),
    .C1(_05217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05218_));
 sky130_fd_sc_hd__a221o_1 _11373_ (.A1(\sha256cu.m_pad_pars.block_512[9][5] ),
    .A2(_05144_),
    .B1(_05147_),
    .B2(\sha256cu.m_pad_pars.block_512[33][5] ),
    .C1(_05218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05219_));
 sky130_fd_sc_hd__or3_1 _11374_ (.A(_05212_),
    .B(_05214_),
    .C(_05219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05220_));
 sky130_fd_sc_hd__a22o_1 _11375_ (.A1(\sha256cu.data_in_padd[21] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00884_));
 sky130_fd_sc_hd__a22o_1 _11376_ (.A1(\sha256cu.m_pad_pars.block_512[13][6] ),
    .A2(_05128_),
    .B1(_05144_),
    .B2(\sha256cu.m_pad_pars.block_512[9][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05221_));
 sky130_fd_sc_hd__a22o_1 _11377_ (.A1(\sha256cu.m_pad_pars.block_512[25][6] ),
    .A2(_05140_),
    .B1(_05141_),
    .B2(\sha256cu.m_pad_pars.block_512[29][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05222_));
 sky130_fd_sc_hd__a221o_1 _11378_ (.A1(\sha256cu.m_pad_pars.block_512[1][6] ),
    .A2(_05135_),
    .B1(_05138_),
    .B2(\sha256cu.m_pad_pars.block_512[17][6] ),
    .C1(_05222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05223_));
 sky130_fd_sc_hd__a22o_1 _11379_ (.A1(\sha256cu.m_pad_pars.block_512[61][6] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05224_));
 sky130_fd_sc_hd__a22o_1 _11380_ (.A1(\sha256cu.m_pad_pars.block_512[53][6] ),
    .A2(_05161_),
    .B1(_05224_),
    .B2(_05024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05225_));
 sky130_fd_sc_hd__a221o_1 _11381_ (.A1(\sha256cu.m_pad_pars.block_512[5][6] ),
    .A2(_05160_),
    .B1(_05165_),
    .B2(\sha256cu.m_pad_pars.block_512[37][6] ),
    .C1(_05225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05226_));
 sky130_fd_sc_hd__a221o_1 _11382_ (.A1(\sha256cu.m_pad_pars.block_512[49][6] ),
    .A2(_05151_),
    .B1(_05158_),
    .B2(\sha256cu.m_pad_pars.block_512[21][6] ),
    .C1(_05226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05227_));
 sky130_fd_sc_hd__a22o_1 _11383_ (.A1(\sha256cu.m_pad_pars.block_512[41][6] ),
    .A2(_05132_),
    .B1(_05147_),
    .B2(\sha256cu.m_pad_pars.block_512[33][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05228_));
 sky130_fd_sc_hd__or3_1 _11384_ (.A(_05223_),
    .B(_05227_),
    .C(_05228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05229_));
 sky130_fd_sc_hd__a211o_1 _11385_ (.A1(\sha256cu.m_pad_pars.block_512[45][6] ),
    .A2(_05126_),
    .B1(_05221_),
    .C1(_05229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05230_));
 sky130_fd_sc_hd__a22o_1 _11386_ (.A1(\sha256cu.data_in_padd[22] ),
    .A2(_04741_),
    .B1(_04742_),
    .B2(_05230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00885_));
 sky130_fd_sc_hd__nor2_1 _11387_ (.A(_04794_),
    .B(_04960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05231_));
 sky130_fd_sc_hd__o22a_1 _11388_ (.A1(_04917_),
    .A2(_05129_),
    .B1(_05231_),
    .B2(\sha256cu.m_pad_pars.block_512[41][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05232_));
 sky130_fd_sc_hd__or2_1 _11389_ (.A(_04704_),
    .B(_05154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05233_));
 sky130_fd_sc_hd__nor2_1 _11390_ (.A(_04824_),
    .B(_04969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05234_));
 sky130_fd_sc_hd__o22a_1 _11391_ (.A1(_01952_),
    .A2(_05233_),
    .B1(_05234_),
    .B2(\sha256cu.m_pad_pars.block_512[53][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05235_));
 sky130_fd_sc_hd__o22a_1 _11392_ (.A1(_04747_),
    .A2(_05154_),
    .B1(_05155_),
    .B2(\sha256cu.m_pad_pars.block_512[21][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05236_));
 sky130_fd_sc_hd__and3b_1 _11393_ (.A_N(_04954_),
    .B(_01956_),
    .C(_04786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05237_));
 sky130_fd_sc_hd__o22a_1 _11394_ (.A1(_04768_),
    .A2(_05154_),
    .B1(_05237_),
    .B2(\sha256cu.m_pad_pars.block_512[5][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05238_));
 sky130_fd_sc_hd__and3_1 _11395_ (.A(_05127_),
    .B(_05152_),
    .C(_05238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05239_));
 sky130_fd_sc_hd__a31o_1 _11396_ (.A1(_01985_),
    .A2(_05152_),
    .A3(_05236_),
    .B1(_05239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05240_));
 sky130_fd_sc_hd__a31o_1 _11397_ (.A1(_05152_),
    .A2(_05149_),
    .A3(_05235_),
    .B1(_05240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05241_));
 sky130_fd_sc_hd__nor2_1 _11398_ (.A(_04960_),
    .B(_05010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05242_));
 sky130_fd_sc_hd__o22a_1 _11399_ (.A1(_04907_),
    .A2(_05129_),
    .B1(_05242_),
    .B2(\sha256cu.m_pad_pars.block_512[25][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05243_));
 sky130_fd_sc_hd__nor2_1 _11400_ (.A(_04787_),
    .B(_04993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05244_));
 sky130_fd_sc_hd__o211a_1 _11401_ (.A1(\sha256cu.m_pad_pars.block_512[1][7] ),
    .A2(_05244_),
    .B1(_05134_),
    .C1(_05127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05245_));
 sky130_fd_sc_hd__nor2_1 _11402_ (.A(_04792_),
    .B(_04969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05246_));
 sky130_fd_sc_hd__o22a_1 _11403_ (.A1(_04819_),
    .A2(_05233_),
    .B1(_05246_),
    .B2(\sha256cu.m_pad_pars.block_512[37][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05247_));
 sky130_fd_sc_hd__or2_2 _11404_ (.A(_01941_),
    .B(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05248_));
 sky130_fd_sc_hd__o21a_1 _11405_ (.A1(_04746_),
    .A2(_05248_),
    .B1(\sha256cu.m_pad_pars.block_512[29][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05249_));
 sky130_fd_sc_hd__a31o_1 _11406_ (.A1(_04699_),
    .A2(_04925_),
    .A3(_04973_),
    .B1(_05249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05250_));
 sky130_fd_sc_hd__and3_1 _11407_ (.A(_01977_),
    .B(_01985_),
    .C(_05250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05251_));
 sky130_fd_sc_hd__a31o_1 _11408_ (.A1(_05125_),
    .A2(_05152_),
    .A3(_05247_),
    .B1(_05251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05252_));
 sky130_fd_sc_hd__a311o_1 _11409_ (.A1(_01985_),
    .A2(_05139_),
    .A3(_05243_),
    .B1(_05245_),
    .C1(_05252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05253_));
 sky130_fd_sc_hd__a311o_1 _11410_ (.A1(_05125_),
    .A2(_05139_),
    .A3(_05232_),
    .B1(_05241_),
    .C1(_05253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05254_));
 sky130_fd_sc_hd__o21a_1 _11411_ (.A1(_04917_),
    .A2(_05248_),
    .B1(\sha256cu.m_pad_pars.block_512[45][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05255_));
 sky130_fd_sc_hd__a31o_1 _11412_ (.A1(_04698_),
    .A2(_04801_),
    .A3(_04973_),
    .B1(_05255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05256_));
 sky130_fd_sc_hd__nor2_1 _11413_ (.A(_04702_),
    .B(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05257_));
 sky130_fd_sc_hd__o22a_1 _11414_ (.A1(_04933_),
    .A2(_05248_),
    .B1(_05257_),
    .B2(\sha256cu.m_pad_pars.block_512[13][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05258_));
 sky130_fd_sc_hd__nor2_1 _11415_ (.A(_04702_),
    .B(_05091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05259_));
 sky130_fd_sc_hd__o22a_1 _11416_ (.A1(_04769_),
    .A2(_05129_),
    .B1(_05259_),
    .B2(\sha256cu.m_pad_pars.block_512[9][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05260_));
 sky130_fd_sc_hd__and3_1 _11417_ (.A(_05127_),
    .B(_05139_),
    .C(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05261_));
 sky130_fd_sc_hd__a31o_1 _11418_ (.A1(_01977_),
    .A2(_05127_),
    .A3(_05258_),
    .B1(_05261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05262_));
 sky130_fd_sc_hd__a31o_1 _11419_ (.A1(_01977_),
    .A2(_05125_),
    .A3(_05256_),
    .B1(_05262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05263_));
 sky130_fd_sc_hd__or2_1 _11420_ (.A(_01940_),
    .B(_01941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05264_));
 sky130_fd_sc_hd__nor2_1 _11421_ (.A(_04807_),
    .B(_05004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05265_));
 sky130_fd_sc_hd__o22a_1 _11422_ (.A1(_05264_),
    .A2(_04907_),
    .B1(_05265_),
    .B2(\sha256cu.m_pad_pars.block_512[17][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05266_));
 sky130_fd_sc_hd__o22a_1 _11423_ (.A1(_05264_),
    .A2(_04913_),
    .B1(_05145_),
    .B2(\sha256cu.m_pad_pars.block_512[33][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05267_));
 sky130_fd_sc_hd__a22o_1 _11424_ (.A1(\sha256cu.m_pad_pars.block_512[61][7] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\sha256cu.m_pad_pars.block_512[57][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05268_));
 sky130_fd_sc_hd__nor2_1 _11425_ (.A(_04824_),
    .B(_05004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05269_));
 sky130_fd_sc_hd__o22a_1 _11426_ (.A1(_01950_),
    .A2(_05136_),
    .B1(_05269_),
    .B2(\sha256cu.m_pad_pars.block_512[49][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05270_));
 sky130_fd_sc_hd__a22o_1 _11427_ (.A1(_01920_),
    .A2(_05268_),
    .B1(_05270_),
    .B2(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05271_));
 sky130_fd_sc_hd__a31o_1 _11428_ (.A1(_05125_),
    .A2(_05134_),
    .A3(_05267_),
    .B1(_05271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05272_));
 sky130_fd_sc_hd__a311o_1 _11429_ (.A1(_01985_),
    .A2(_05134_),
    .A3(_05266_),
    .B1(_05272_),
    .C1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05273_));
 sky130_fd_sc_hd__or3_1 _11430_ (.A(_05254_),
    .B(_05263_),
    .C(_05273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05274_));
 sky130_fd_sc_hd__o211a_1 _11431_ (.A1(\sha256cu.data_in_padd[23] ),
    .A2(_04840_),
    .B1(_05274_),
    .C1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00886_));
 sky130_fd_sc_hd__nor2_2 _11432_ (.A(_04701_),
    .B(_05129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05275_));
 sky130_fd_sc_hd__nor2_1 _11433_ (.A(_04924_),
    .B(_05275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05276_));
 sky130_fd_sc_hd__nor2b_2 _11434_ (.A(\sha256cu.m_pad_pars.add_out0[5] ),
    .B_N(\sha256cu.m_pad_pars.add_out0[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05277_));
 sky130_fd_sc_hd__nor2b_2 _11435_ (.A(\sha256cu.m_pad_pars.add_out0[2] ),
    .B_N(\sha256cu.m_pad_pars.add_out0[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05278_));
 sky130_fd_sc_hd__o211a_2 _11436_ (.A1(_04907_),
    .A2(_05276_),
    .B1(_05277_),
    .C1(_05278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05279_));
 sky130_fd_sc_hd__and3_2 _11437_ (.A(\sha256cu.m_pad_pars.add_out0[5] ),
    .B(\sha256cu.m_pad_pars.add_out0[4] ),
    .C(_05278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05280_));
 sky130_fd_sc_hd__a22o_1 _11438_ (.A1(\sha256cu.m_pad_pars.block_512[60][0] ),
    .A2(_01998_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05281_));
 sky130_fd_sc_hd__nor2_1 _11439_ (.A(_04807_),
    .B(_05136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05282_));
 sky130_fd_sc_hd__a31o_1 _11440_ (.A1(_01944_),
    .A2(_04699_),
    .A3(_04777_),
    .B1(_05282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05283_));
 sky130_fd_sc_hd__inv_1 _11441_ (.A(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05284_));
 sky130_fd_sc_hd__and3_2 _11442_ (.A(_01935_),
    .B(_05277_),
    .C(_05284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05285_));
 sky130_fd_sc_hd__o22a_1 _11443_ (.A1(_04808_),
    .A2(_04819_),
    .B1(_04824_),
    .B2(_05264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05286_));
 sky130_fd_sc_hd__and3_1 _11444_ (.A(\sha256cu.m_pad_pars.add_out0[5] ),
    .B(\sha256cu.m_pad_pars.add_out0[4] ),
    .C(_01935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05287_));
 sky130_fd_sc_hd__o21a_2 _11445_ (.A1(_04705_),
    .A2(_05286_),
    .B1(_05287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05288_));
 sky130_fd_sc_hd__a22o_1 _11446_ (.A1(\sha256cu.m_pad_pars.block_512[16][0] ),
    .A2(_05285_),
    .B1(_05288_),
    .B2(\sha256cu.m_pad_pars.block_512[48][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05289_));
 sky130_fd_sc_hd__a221o_1 _11447_ (.A1(\sha256cu.m_pad_pars.block_512[24][0] ),
    .A2(_05279_),
    .B1(_05281_),
    .B2(_01921_),
    .C1(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05290_));
 sky130_fd_sc_hd__nor2_1 _11448_ (.A(_04701_),
    .B(_05154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05291_));
 sky130_fd_sc_hd__nor2_1 _11449_ (.A(_04760_),
    .B(_05291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05292_));
 sky130_fd_sc_hd__and2b_2 _11450_ (.A_N(\sha256cu.m_pad_pars.add_out0[3] ),
    .B(\sha256cu.m_pad_pars.add_out0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05293_));
 sky130_fd_sc_hd__o211a_2 _11451_ (.A1(_04907_),
    .A2(_05292_),
    .B1(_05293_),
    .C1(_05277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05294_));
 sky130_fd_sc_hd__o21a_1 _11452_ (.A1(_04701_),
    .A2(_05248_),
    .B1(_04751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05295_));
 sky130_fd_sc_hd__o211a_2 _11453_ (.A1(_04746_),
    .A2(_05295_),
    .B1(_05277_),
    .C1(_01992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05296_));
 sky130_fd_sc_hd__nor2b_2 _11454_ (.A(\sha256cu.m_pad_pars.add_out0[4] ),
    .B_N(\sha256cu.m_pad_pars.add_out0[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05297_));
 sky130_fd_sc_hd__o211a_2 _11455_ (.A1(_04912_),
    .A2(_05295_),
    .B1(_05297_),
    .C1(_01992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05298_));
 sky130_fd_sc_hd__o211a_2 _11456_ (.A1(_04769_),
    .A2(_05295_),
    .B1(_01936_),
    .C1(_01992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05299_));
 sky130_fd_sc_hd__a22o_1 _11457_ (.A1(\sha256cu.m_pad_pars.block_512[44][0] ),
    .A2(_05298_),
    .B1(_05299_),
    .B2(\sha256cu.m_pad_pars.block_512[12][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05300_));
 sky130_fd_sc_hd__a221o_1 _11458_ (.A1(\sha256cu.m_pad_pars.block_512[20][0] ),
    .A2(_05294_),
    .B1(_05296_),
    .B2(\sha256cu.m_pad_pars.block_512[28][0] ),
    .C1(_05300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05301_));
 sky130_fd_sc_hd__nor2_1 _11459_ (.A(_04794_),
    .B(_05154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05302_));
 sky130_fd_sc_hd__a21oi_1 _11460_ (.A1(_04760_),
    .A2(_04801_),
    .B1(_05302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05303_));
 sky130_fd_sc_hd__and3_2 _11461_ (.A(_05293_),
    .B(_05297_),
    .C(_05303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05304_));
 sky130_fd_sc_hd__o21a_1 _11462_ (.A1(_04792_),
    .A2(_05136_),
    .B1(_04909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05305_));
 sky130_fd_sc_hd__and3_2 _11463_ (.A(_01935_),
    .B(_05297_),
    .C(_05305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05306_));
 sky130_fd_sc_hd__or3_1 _11464_ (.A(_04703_),
    .B(_04824_),
    .C(_05154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05307_));
 sky130_fd_sc_hd__o21ai_1 _11465_ (.A1(_01952_),
    .A2(_04761_),
    .B1(_05307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05308_));
 sky130_fd_sc_hd__inv_1 _11466_ (.A(_05308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05309_));
 sky130_fd_sc_hd__and4_2 _11467_ (.A(\sha256cu.m_pad_pars.add_out0[5] ),
    .B(\sha256cu.m_pad_pars.add_out0[4] ),
    .C(_05293_),
    .D(_05309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05310_));
 sky130_fd_sc_hd__a22o_1 _11468_ (.A1(\sha256cu.m_pad_pars.block_512[32][0] ),
    .A2(_05306_),
    .B1(_05310_),
    .B2(\sha256cu.m_pad_pars.block_512[52][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05311_));
 sky130_fd_sc_hd__o32a_1 _11469_ (.A1(_04701_),
    .A2(_04768_),
    .A3(_05154_),
    .B1(_01943_),
    .B2(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05312_));
 sky130_fd_sc_hd__and3_2 _11470_ (.A(_01936_),
    .B(_05293_),
    .C(_05312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05313_));
 sky130_fd_sc_hd__a21oi_4 _11471_ (.A1(_01942_),
    .A2(_04775_),
    .B1(_01937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05314_));
 sky130_fd_sc_hd__nand2_1 _11472_ (.A(_01936_),
    .B(_05278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05315_));
 sky130_fd_sc_hd__nor2_1 _11473_ (.A(\sha256cu.m_pad_pars.add_512_block[6] ),
    .B(_04770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05316_));
 sky130_fd_sc_hd__o21a_1 _11474_ (.A1(_05275_),
    .A2(_05316_),
    .B1(_04786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05317_));
 sky130_fd_sc_hd__nor2_4 _11475_ (.A(_05315_),
    .B(_05317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05318_));
 sky130_fd_sc_hd__o21a_1 _11476_ (.A1(_05275_),
    .A2(_05316_),
    .B1(_04801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05319_));
 sky130_fd_sc_hd__and3b_2 _11477_ (.A_N(_05319_),
    .B(_05297_),
    .C(_05278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05320_));
 sky130_fd_sc_hd__a22o_1 _11478_ (.A1(\sha256cu.m_pad_pars.block_512[8][0] ),
    .A2(_05318_),
    .B1(_05320_),
    .B2(\sha256cu.m_pad_pars.block_512[40][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05321_));
 sky130_fd_sc_hd__a221o_1 _11479_ (.A1(\sha256cu.m_pad_pars.block_512[4][0] ),
    .A2(_05313_),
    .B1(_05314_),
    .B2(\sha256cu.m_pad_pars.block_512[0][0] ),
    .C1(_05321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05322_));
 sky130_fd_sc_hd__a211o_1 _11480_ (.A1(\sha256cu.m_pad_pars.block_512[36][0] ),
    .A2(_05304_),
    .B1(_05311_),
    .C1(_05322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05323_));
 sky130_fd_sc_hd__or3_2 _11481_ (.A(_05290_),
    .B(_05301_),
    .C(_05323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05324_));
 sky130_fd_sc_hd__a22o_1 _11482_ (.A1(\sha256cu.data_in_padd[24] ),
    .A2(_01980_),
    .B1(_01987_),
    .B2(_05324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00887_));
 sky130_fd_sc_hd__a22o_1 _11483_ (.A1(\sha256cu.m_pad_pars.block_512[60][1] ),
    .A2(_01998_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05325_));
 sky130_fd_sc_hd__a22o_1 _11484_ (.A1(\sha256cu.m_pad_pars.block_512[36][1] ),
    .A2(_05304_),
    .B1(_05325_),
    .B2(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05326_));
 sky130_fd_sc_hd__a221o_1 _11485_ (.A1(\sha256cu.m_pad_pars.block_512[8][1] ),
    .A2(_05318_),
    .B1(_05285_),
    .B2(\sha256cu.m_pad_pars.block_512[16][1] ),
    .C1(_05326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05327_));
 sky130_fd_sc_hd__a22o_1 _11486_ (.A1(\sha256cu.m_pad_pars.block_512[24][1] ),
    .A2(_05279_),
    .B1(_05294_),
    .B2(\sha256cu.m_pad_pars.block_512[20][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05328_));
 sky130_fd_sc_hd__a22o_1 _11487_ (.A1(\sha256cu.m_pad_pars.block_512[44][1] ),
    .A2(_05298_),
    .B1(_05296_),
    .B2(\sha256cu.m_pad_pars.block_512[28][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05329_));
 sky130_fd_sc_hd__a221o_1 _11488_ (.A1(\sha256cu.m_pad_pars.block_512[32][1] ),
    .A2(_05306_),
    .B1(_05310_),
    .B2(\sha256cu.m_pad_pars.block_512[52][1] ),
    .C1(_05329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05330_));
 sky130_fd_sc_hd__a22o_1 _11489_ (.A1(\sha256cu.m_pad_pars.block_512[4][1] ),
    .A2(_05313_),
    .B1(_05288_),
    .B2(\sha256cu.m_pad_pars.block_512[48][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05331_));
 sky130_fd_sc_hd__a221o_1 _11490_ (.A1(\sha256cu.m_pad_pars.block_512[40][1] ),
    .A2(_05320_),
    .B1(_05299_),
    .B2(\sha256cu.m_pad_pars.block_512[12][1] ),
    .C1(_05331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05332_));
 sky130_fd_sc_hd__or4_1 _11491_ (.A(_05327_),
    .B(_05328_),
    .C(_05330_),
    .D(_05332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05333_));
 sky130_fd_sc_hd__a211o_1 _11492_ (.A1(\sha256cu.m_pad_pars.block_512[0][1] ),
    .A2(_05314_),
    .B1(_05333_),
    .C1(_01971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05334_));
 sky130_fd_sc_hd__clkbuf_4 _11493_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05335_));
 sky130_fd_sc_hd__o211a_1 _11494_ (.A1(\sha256cu.data_in_padd[25] ),
    .A2(_04840_),
    .B1(_05334_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00888_));
 sky130_fd_sc_hd__a22o_1 _11495_ (.A1(\sha256cu.m_pad_pars.block_512[24][2] ),
    .A2(_05279_),
    .B1(_05298_),
    .B2(\sha256cu.m_pad_pars.block_512[44][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05336_));
 sky130_fd_sc_hd__a221o_1 _11496_ (.A1(\sha256cu.m_pad_pars.block_512[32][2] ),
    .A2(_05306_),
    .B1(_05318_),
    .B2(\sha256cu.m_pad_pars.block_512[8][2] ),
    .C1(_05336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05337_));
 sky130_fd_sc_hd__a22o_1 _11497_ (.A1(\sha256cu.m_pad_pars.block_512[4][2] ),
    .A2(_05313_),
    .B1(_05320_),
    .B2(\sha256cu.m_pad_pars.block_512[40][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05338_));
 sky130_fd_sc_hd__a221o_1 _11498_ (.A1(\sha256cu.m_pad_pars.block_512[12][2] ),
    .A2(_05299_),
    .B1(_05304_),
    .B2(\sha256cu.m_pad_pars.block_512[36][2] ),
    .C1(_05338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05339_));
 sky130_fd_sc_hd__a22o_1 _11499_ (.A1(\sha256cu.m_pad_pars.block_512[20][2] ),
    .A2(_05294_),
    .B1(_05285_),
    .B2(\sha256cu.m_pad_pars.block_512[16][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05340_));
 sky130_fd_sc_hd__a22o_1 _11500_ (.A1(\sha256cu.m_pad_pars.block_512[60][2] ),
    .A2(_01998_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05341_));
 sky130_fd_sc_hd__a22o_1 _11501_ (.A1(\sha256cu.m_pad_pars.block_512[28][2] ),
    .A2(_05296_),
    .B1(_05341_),
    .B2(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05342_));
 sky130_fd_sc_hd__a221o_1 _11502_ (.A1(\sha256cu.m_pad_pars.block_512[52][2] ),
    .A2(_05310_),
    .B1(_05288_),
    .B2(\sha256cu.m_pad_pars.block_512[48][2] ),
    .C1(_05342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05343_));
 sky130_fd_sc_hd__a211o_1 _11503_ (.A1(\sha256cu.m_pad_pars.block_512[0][2] ),
    .A2(_05314_),
    .B1(_05340_),
    .C1(_05343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05344_));
 sky130_fd_sc_hd__or3_2 _11504_ (.A(_05337_),
    .B(_05339_),
    .C(_05344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05345_));
 sky130_fd_sc_hd__a22o_1 _11505_ (.A1(\sha256cu.data_in_padd[26] ),
    .A2(_01980_),
    .B1(_01987_),
    .B2(_05345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00889_));
 sky130_fd_sc_hd__a22o_1 _11506_ (.A1(\sha256cu.m_pad_pars.block_512[24][3] ),
    .A2(_05279_),
    .B1(_05298_),
    .B2(\sha256cu.m_pad_pars.block_512[44][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05346_));
 sky130_fd_sc_hd__a221o_1 _11507_ (.A1(\sha256cu.m_pad_pars.block_512[32][3] ),
    .A2(_05306_),
    .B1(_05318_),
    .B2(\sha256cu.m_pad_pars.block_512[8][3] ),
    .C1(_05346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05347_));
 sky130_fd_sc_hd__a22o_1 _11508_ (.A1(\sha256cu.m_pad_pars.block_512[4][3] ),
    .A2(_05313_),
    .B1(_05320_),
    .B2(\sha256cu.m_pad_pars.block_512[40][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05348_));
 sky130_fd_sc_hd__a221o_1 _11509_ (.A1(\sha256cu.m_pad_pars.block_512[12][3] ),
    .A2(_05299_),
    .B1(_05304_),
    .B2(\sha256cu.m_pad_pars.block_512[36][3] ),
    .C1(_05348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05349_));
 sky130_fd_sc_hd__a22o_1 _11510_ (.A1(\sha256cu.m_pad_pars.block_512[20][3] ),
    .A2(_05294_),
    .B1(_05285_),
    .B2(\sha256cu.m_pad_pars.block_512[16][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05350_));
 sky130_fd_sc_hd__a22o_1 _11511_ (.A1(\sha256cu.m_pad_pars.block_512[60][3] ),
    .A2(_01998_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05351_));
 sky130_fd_sc_hd__a22o_1 _11512_ (.A1(\sha256cu.m_pad_pars.block_512[28][3] ),
    .A2(_05296_),
    .B1(_05351_),
    .B2(_01921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05352_));
 sky130_fd_sc_hd__a221o_1 _11513_ (.A1(\sha256cu.m_pad_pars.block_512[52][3] ),
    .A2(_05310_),
    .B1(_05288_),
    .B2(\sha256cu.m_pad_pars.block_512[48][3] ),
    .C1(_05352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05353_));
 sky130_fd_sc_hd__a211o_1 _11514_ (.A1(\sha256cu.m_pad_pars.block_512[0][3] ),
    .A2(_05314_),
    .B1(_05350_),
    .C1(_05353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05354_));
 sky130_fd_sc_hd__or3_2 _11515_ (.A(_05347_),
    .B(_05349_),
    .C(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05355_));
 sky130_fd_sc_hd__a22o_1 _11516_ (.A1(\sha256cu.data_in_padd[27] ),
    .A2(_01980_),
    .B1(_01987_),
    .B2(_05355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00890_));
 sky130_fd_sc_hd__a22o_1 _11517_ (.A1(\sha256cu.m_pad_pars.block_512[24][4] ),
    .A2(_05279_),
    .B1(_05313_),
    .B2(\sha256cu.m_pad_pars.block_512[4][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05356_));
 sky130_fd_sc_hd__a221o_1 _11518_ (.A1(\sha256cu.m_pad_pars.block_512[32][4] ),
    .A2(_05306_),
    .B1(_05318_),
    .B2(\sha256cu.m_pad_pars.block_512[8][4] ),
    .C1(_05356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05357_));
 sky130_fd_sc_hd__a22o_1 _11519_ (.A1(\sha256cu.m_pad_pars.block_512[44][4] ),
    .A2(_05298_),
    .B1(_05320_),
    .B2(\sha256cu.m_pad_pars.block_512[40][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05358_));
 sky130_fd_sc_hd__a221o_1 _11520_ (.A1(\sha256cu.m_pad_pars.block_512[12][4] ),
    .A2(_05299_),
    .B1(_05304_),
    .B2(\sha256cu.m_pad_pars.block_512[36][4] ),
    .C1(_05358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05359_));
 sky130_fd_sc_hd__a22o_1 _11521_ (.A1(\sha256cu.m_pad_pars.block_512[20][4] ),
    .A2(_05294_),
    .B1(_05285_),
    .B2(\sha256cu.m_pad_pars.block_512[16][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05360_));
 sky130_fd_sc_hd__a22o_1 _11522_ (.A1(\sha256cu.m_pad_pars.block_512[60][4] ),
    .A2(_01998_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05361_));
 sky130_fd_sc_hd__a22o_1 _11523_ (.A1(\sha256cu.m_pad_pars.block_512[28][4] ),
    .A2(_05296_),
    .B1(_05361_),
    .B2(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05362_));
 sky130_fd_sc_hd__a221o_1 _11524_ (.A1(\sha256cu.m_pad_pars.block_512[52][4] ),
    .A2(_05310_),
    .B1(_05288_),
    .B2(\sha256cu.m_pad_pars.block_512[48][4] ),
    .C1(_05362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05363_));
 sky130_fd_sc_hd__a211o_1 _11525_ (.A1(\sha256cu.m_pad_pars.block_512[0][4] ),
    .A2(_05314_),
    .B1(_05360_),
    .C1(_05363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05364_));
 sky130_fd_sc_hd__or3_2 _11526_ (.A(_05357_),
    .B(_05359_),
    .C(_05364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05365_));
 sky130_fd_sc_hd__a22o_1 _11527_ (.A1(\sha256cu.data_in_padd[28] ),
    .A2(_01980_),
    .B1(_01987_),
    .B2(_05365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00891_));
 sky130_fd_sc_hd__a22o_1 _11528_ (.A1(\sha256cu.m_pad_pars.block_512[24][5] ),
    .A2(_05279_),
    .B1(_05304_),
    .B2(\sha256cu.m_pad_pars.block_512[36][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05366_));
 sky130_fd_sc_hd__a221o_1 _11529_ (.A1(\sha256cu.m_pad_pars.block_512[32][5] ),
    .A2(_05306_),
    .B1(_05318_),
    .B2(\sha256cu.m_pad_pars.block_512[8][5] ),
    .C1(_05366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05367_));
 sky130_fd_sc_hd__a22o_1 _11530_ (.A1(\sha256cu.m_pad_pars.block_512[4][5] ),
    .A2(_05313_),
    .B1(_05299_),
    .B2(\sha256cu.m_pad_pars.block_512[12][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05368_));
 sky130_fd_sc_hd__a221o_1 _11531_ (.A1(\sha256cu.m_pad_pars.block_512[44][5] ),
    .A2(_05298_),
    .B1(_05320_),
    .B2(\sha256cu.m_pad_pars.block_512[40][5] ),
    .C1(_05368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05369_));
 sky130_fd_sc_hd__a22o_1 _11532_ (.A1(\sha256cu.m_pad_pars.block_512[16][5] ),
    .A2(_05285_),
    .B1(_05296_),
    .B2(\sha256cu.m_pad_pars.block_512[28][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05370_));
 sky130_fd_sc_hd__a22o_1 _11533_ (.A1(\sha256cu.m_pad_pars.block_512[60][5] ),
    .A2(_01998_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05371_));
 sky130_fd_sc_hd__a22o_1 _11534_ (.A1(\sha256cu.m_pad_pars.block_512[52][5] ),
    .A2(_05310_),
    .B1(_05371_),
    .B2(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05372_));
 sky130_fd_sc_hd__a221o_1 _11535_ (.A1(\sha256cu.m_pad_pars.block_512[20][5] ),
    .A2(_05294_),
    .B1(_05288_),
    .B2(\sha256cu.m_pad_pars.block_512[48][5] ),
    .C1(_05372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05373_));
 sky130_fd_sc_hd__a211o_1 _11536_ (.A1(\sha256cu.m_pad_pars.block_512[0][5] ),
    .A2(_05314_),
    .B1(_05370_),
    .C1(_05373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05374_));
 sky130_fd_sc_hd__or3_2 _11537_ (.A(_05367_),
    .B(_05369_),
    .C(_05374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05375_));
 sky130_fd_sc_hd__a22o_1 _11538_ (.A1(\sha256cu.data_in_padd[29] ),
    .A2(_01980_),
    .B1(_01987_),
    .B2(_05375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00892_));
 sky130_fd_sc_hd__a22o_1 _11539_ (.A1(\sha256cu.m_pad_pars.block_512[8][6] ),
    .A2(_05318_),
    .B1(_05299_),
    .B2(\sha256cu.m_pad_pars.block_512[12][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05376_));
 sky130_fd_sc_hd__a221o_1 _11540_ (.A1(\sha256cu.m_pad_pars.block_512[32][6] ),
    .A2(_05306_),
    .B1(_05320_),
    .B2(\sha256cu.m_pad_pars.block_512[40][6] ),
    .C1(_05376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05377_));
 sky130_fd_sc_hd__a22o_1 _11541_ (.A1(\sha256cu.m_pad_pars.block_512[24][6] ),
    .A2(_05279_),
    .B1(_05313_),
    .B2(\sha256cu.m_pad_pars.block_512[4][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05378_));
 sky130_fd_sc_hd__a221o_1 _11542_ (.A1(\sha256cu.m_pad_pars.block_512[44][6] ),
    .A2(_05298_),
    .B1(_05304_),
    .B2(\sha256cu.m_pad_pars.block_512[36][6] ),
    .C1(_05378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05379_));
 sky130_fd_sc_hd__a22o_1 _11543_ (.A1(\sha256cu.m_pad_pars.block_512[16][6] ),
    .A2(_05285_),
    .B1(_05288_),
    .B2(\sha256cu.m_pad_pars.block_512[48][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05380_));
 sky130_fd_sc_hd__a22o_1 _11544_ (.A1(\sha256cu.m_pad_pars.block_512[60][6] ),
    .A2(_01998_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05381_));
 sky130_fd_sc_hd__a22o_1 _11545_ (.A1(\sha256cu.m_pad_pars.block_512[28][6] ),
    .A2(_05296_),
    .B1(_05381_),
    .B2(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05382_));
 sky130_fd_sc_hd__a221o_1 _11546_ (.A1(\sha256cu.m_pad_pars.block_512[20][6] ),
    .A2(_05294_),
    .B1(_05314_),
    .B2(\sha256cu.m_pad_pars.block_512[0][6] ),
    .C1(_05382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05383_));
 sky130_fd_sc_hd__a211o_1 _11547_ (.A1(\sha256cu.m_pad_pars.block_512[52][6] ),
    .A2(_05310_),
    .B1(_05380_),
    .C1(_05383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05384_));
 sky130_fd_sc_hd__or3_2 _11548_ (.A(_05377_),
    .B(_05379_),
    .C(_05384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05385_));
 sky130_fd_sc_hd__a22o_1 _11549_ (.A1(\sha256cu.data_in_padd[30] ),
    .A2(_01980_),
    .B1(_01987_),
    .B2(_05385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00893_));
 sky130_fd_sc_hd__inv_2 _11550_ (.A(_05314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05386_));
 sky130_fd_sc_hd__nor2_1 _11551_ (.A(_05010_),
    .B(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05387_));
 sky130_fd_sc_hd__o22a_1 _11552_ (.A1(_04907_),
    .A2(_04751_),
    .B1(_05387_),
    .B2(\sha256cu.m_pad_pars.block_512[28][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05388_));
 sky130_fd_sc_hd__nor2_1 _11553_ (.A(_04794_),
    .B(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05389_));
 sky130_fd_sc_hd__o22a_1 _11554_ (.A1(_04751_),
    .A2(_04917_),
    .B1(_05389_),
    .B2(\sha256cu.m_pad_pars.block_512[44][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05390_));
 sky130_fd_sc_hd__a22o_1 _11555_ (.A1(_05277_),
    .A2(_05388_),
    .B1(_05390_),
    .B2(_05297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05391_));
 sky130_fd_sc_hd__and2_1 _11556_ (.A(_01992_),
    .B(_05391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05392_));
 sky130_fd_sc_hd__nor2_1 _11557_ (.A(_04792_),
    .B(_05136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05393_));
 sky130_fd_sc_hd__o21a_1 _11558_ (.A1(\sha256cu.m_pad_pars.block_512[32][7] ),
    .A2(_05393_),
    .B1(_04909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05394_));
 sky130_fd_sc_hd__nor2_1 _11559_ (.A(_04807_),
    .B(_05233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05395_));
 sky130_fd_sc_hd__o22a_1 _11560_ (.A1(_04747_),
    .A2(_04815_),
    .B1(_05395_),
    .B2(\sha256cu.m_pad_pars.block_512[20][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05396_));
 sky130_fd_sc_hd__and3_1 _11561_ (.A(_05277_),
    .B(_05293_),
    .C(_05396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05397_));
 sky130_fd_sc_hd__a31o_1 _11562_ (.A1(_01935_),
    .A2(_05297_),
    .A3(_05394_),
    .B1(_05397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05398_));
 sky130_fd_sc_hd__a21oi_1 _11563_ (.A1(_04801_),
    .A2(_05275_),
    .B1(\sha256cu.m_pad_pars.block_512[40][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05399_));
 sky130_fd_sc_hd__a21oi_1 _11564_ (.A1(_04801_),
    .A2(_05316_),
    .B1(_05399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05400_));
 sky130_fd_sc_hd__o22a_1 _11565_ (.A1(_04815_),
    .A2(_04913_),
    .B1(_05302_),
    .B2(\sha256cu.m_pad_pars.block_512[36][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05401_));
 sky130_fd_sc_hd__and3_1 _11566_ (.A(_05293_),
    .B(_05297_),
    .C(_05401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05402_));
 sky130_fd_sc_hd__a31o_1 _11567_ (.A1(_05278_),
    .A2(_05297_),
    .A3(_05400_),
    .B1(_05402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05403_));
 sky130_fd_sc_hd__a21oi_1 _11568_ (.A1(_04908_),
    .A2(_05275_),
    .B1(\sha256cu.m_pad_pars.block_512[24][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05404_));
 sky130_fd_sc_hd__a21oi_1 _11569_ (.A1(_04908_),
    .A2(_04924_),
    .B1(_05404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05405_));
 sky130_fd_sc_hd__and3b_1 _11570_ (.A_N(_05248_),
    .B(_04698_),
    .C(_04786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05406_));
 sky130_fd_sc_hd__o22a_1 _11571_ (.A1(_04751_),
    .A2(_04769_),
    .B1(_05406_),
    .B2(\sha256cu.m_pad_pars.block_512[12][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05407_));
 sky130_fd_sc_hd__and3_1 _11572_ (.A(_01936_),
    .B(_01992_),
    .C(_05407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05408_));
 sky130_fd_sc_hd__a31o_1 _11573_ (.A1(_05278_),
    .A2(_05277_),
    .A3(_05405_),
    .B1(_05408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05409_));
 sky130_fd_sc_hd__a21oi_1 _11574_ (.A1(_04786_),
    .A2(_05291_),
    .B1(\sha256cu.m_pad_pars.block_512[4][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05410_));
 sky130_fd_sc_hd__nor2_1 _11575_ (.A(_04762_),
    .B(_05410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05411_));
 sky130_fd_sc_hd__and3_1 _11576_ (.A(_01936_),
    .B(_05293_),
    .C(_05411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05412_));
 sky130_fd_sc_hd__o22a_1 _11577_ (.A1(_04769_),
    .A2(_04808_),
    .B1(_05282_),
    .B2(\sha256cu.m_pad_pars.block_512[16][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05413_));
 sky130_fd_sc_hd__inv_1 _11578_ (.A(\sha256cu.m_pad_pars.block_512[52][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05414_));
 sky130_fd_sc_hd__o2bb2a_1 _11579_ (.A1_N(_05414_),
    .A2_N(_05307_),
    .B1(_04761_),
    .B2(_01952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05415_));
 sky130_fd_sc_hd__inv_2 _11580_ (.A(_01937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05416_));
 sky130_fd_sc_hd__a41o_1 _11581_ (.A1(\sha256cu.m_pad_pars.add_out0[5] ),
    .A2(\sha256cu.m_pad_pars.add_out0[4] ),
    .A3(_05293_),
    .A4(_05415_),
    .B1(_05416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05417_));
 sky130_fd_sc_hd__a31o_1 _11582_ (.A1(_01935_),
    .A2(_05277_),
    .A3(_05413_),
    .B1(_05417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05418_));
 sky130_fd_sc_hd__a22o_1 _11583_ (.A1(\sha256cu.m_pad_pars.block_512[60][7] ),
    .A2(_01997_),
    .B1(_05280_),
    .B2(\sha256cu.m_pad_pars.block_512[56][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05419_));
 sky130_fd_sc_hd__nor2_1 _11584_ (.A(_04824_),
    .B(_05136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05420_));
 sky130_fd_sc_hd__o22a_1 _11585_ (.A1(_04808_),
    .A2(_04912_),
    .B1(_05420_),
    .B2(\sha256cu.m_pad_pars.block_512[48][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05421_));
 sky130_fd_sc_hd__a22o_1 _11586_ (.A1(_01920_),
    .A2(_05419_),
    .B1(_05421_),
    .B2(_05287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05422_));
 sky130_fd_sc_hd__a21oi_1 _11587_ (.A1(_04786_),
    .A2(_05275_),
    .B1(\sha256cu.m_pad_pars.block_512[8][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05423_));
 sky130_fd_sc_hd__a21oi_1 _11588_ (.A1(_04786_),
    .A2(_04924_),
    .B1(_05423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05424_));
 sky130_fd_sc_hd__or2b_1 _11589_ (.A(_05315_),
    .B_N(_05424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05425_));
 sky130_fd_sc_hd__or4b_1 _11590_ (.A(_05412_),
    .B(_05418_),
    .C(_05422_),
    .D_N(_05425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05426_));
 sky130_fd_sc_hd__or4_1 _11591_ (.A(_05398_),
    .B(_05403_),
    .C(_05409_),
    .D(_05426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05427_));
 sky130_fd_sc_hd__o22a_1 _11592_ (.A1(\sha256cu.m_pad_pars.block_512[0][7] ),
    .A2(_05386_),
    .B1(_05392_),
    .B2(_05427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05428_));
 sky130_fd_sc_hd__a22o_1 _11593_ (.A1(\sha256cu.data_in_padd[31] ),
    .A2(_01980_),
    .B1(_01987_),
    .B2(_05428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00894_));
 sky130_fd_sc_hd__and2_1 _11594_ (.A(_03288_),
    .B(_02009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_1 _11595_ (.A(_05429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00895_));
 sky130_fd_sc_hd__a21oi_1 _11596_ (.A1(_04698_),
    .A2(_04705_),
    .B1(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00897_));
 sky130_fd_sc_hd__clkbuf_4 _11597_ (.A(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05430_));
 sky130_fd_sc_hd__a21o_1 _11598_ (.A1(\sha256cu.msg_scheduler.counter_iteration[4] ),
    .A2(_01565_),
    .B1(_04716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05431_));
 sky130_fd_sc_hd__nor4_4 _11599_ (.A(\sha256cu.flag_0_15 ),
    .B(\sha256cu.msg_scheduler.counter_iteration[6] ),
    .C(\sha256cu.msg_scheduler.counter_iteration[5] ),
    .D(_05431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05432_));
 sky130_fd_sc_hd__clkbuf_4 _11600_ (.A(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05433_));
 sky130_fd_sc_hd__nand2_1 _11601_ (.A(\sha256cu.msg_scheduler.mreg_9[0] ),
    .B(\sha256cu.msg_scheduler.mreg_0[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05434_));
 sky130_fd_sc_hd__or2_1 _11602_ (.A(\sha256cu.msg_scheduler.mreg_9[0] ),
    .B(\sha256cu.msg_scheduler.mreg_0[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05435_));
 sky130_fd_sc_hd__nand2_1 _11603_ (.A(_05434_),
    .B(_05435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05436_));
 sky130_fd_sc_hd__xnor2_1 _11604_ (.A(\sha256cu.msg_scheduler.mreg_1[7] ),
    .B(\sha256cu.msg_scheduler.mreg_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05437_));
 sky130_fd_sc_hd__xnor2_1 _11605_ (.A(\sha256cu.msg_scheduler.mreg_1[18] ),
    .B(_05437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05438_));
 sky130_fd_sc_hd__xnor2_1 _11606_ (.A(_05436_),
    .B(_05438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05439_));
 sky130_fd_sc_hd__xnor2_1 _11607_ (.A(\sha256cu.msg_scheduler.mreg_14[17] ),
    .B(\sha256cu.msg_scheduler.mreg_14[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05440_));
 sky130_fd_sc_hd__xnor2_1 _11608_ (.A(\sha256cu.msg_scheduler.mreg_14[19] ),
    .B(_05440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05441_));
 sky130_fd_sc_hd__or4_4 _11609_ (.A(\sha256cu.flag_0_15 ),
    .B(\sha256cu.msg_scheduler.counter_iteration[6] ),
    .C(\sha256cu.msg_scheduler.counter_iteration[5] ),
    .D(_05431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05442_));
 sky130_fd_sc_hd__o21a_1 _11610_ (.A1(_05439_),
    .A2(_05441_),
    .B1(_05442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05443_));
 sky130_fd_sc_hd__nand2_1 _11611_ (.A(_05439_),
    .B(_05441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05444_));
 sky130_fd_sc_hd__clkbuf_4 _11612_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05445_));
 sky130_fd_sc_hd__a221o_1 _11613_ (.A1(\sha256cu.data_in_padd[0] ),
    .A2(_05433_),
    .B1(_05443_),
    .B2(_05444_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05446_));
 sky130_fd_sc_hd__o211a_1 _11614_ (.A1(\sha256cu.iter_processing.w[0] ),
    .A2(_05430_),
    .B1(_05446_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00898_));
 sky130_fd_sc_hd__clkbuf_4 _11615_ (.A(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05447_));
 sky130_fd_sc_hd__buf_2 _11616_ (.A(_05447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05448_));
 sky130_fd_sc_hd__nand2_1 _11617_ (.A(\sha256cu.msg_scheduler.mreg_9[1] ),
    .B(\sha256cu.msg_scheduler.mreg_0[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05449_));
 sky130_fd_sc_hd__or2_1 _11618_ (.A(\sha256cu.msg_scheduler.mreg_9[1] ),
    .B(\sha256cu.msg_scheduler.mreg_0[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_1 _11619_ (.A(_05449_),
    .B(_05450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05451_));
 sky130_fd_sc_hd__xnor2_1 _11620_ (.A(\sha256cu.msg_scheduler.mreg_1[8] ),
    .B(\sha256cu.msg_scheduler.mreg_1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05452_));
 sky130_fd_sc_hd__xnor2_2 _11621_ (.A(\sha256cu.msg_scheduler.mreg_1[19] ),
    .B(_05452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05453_));
 sky130_fd_sc_hd__xor2_2 _11622_ (.A(_05451_),
    .B(_05453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05454_));
 sky130_fd_sc_hd__a21boi_1 _11623_ (.A1(_05435_),
    .A2(_05438_),
    .B1_N(_05434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05455_));
 sky130_fd_sc_hd__xor2_2 _11624_ (.A(_05454_),
    .B(_05455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05456_));
 sky130_fd_sc_hd__xnor2_1 _11625_ (.A(\sha256cu.msg_scheduler.mreg_14[18] ),
    .B(\sha256cu.msg_scheduler.mreg_14[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05457_));
 sky130_fd_sc_hd__xnor2_1 _11626_ (.A(\sha256cu.msg_scheduler.mreg_14[20] ),
    .B(_05457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05458_));
 sky130_fd_sc_hd__xnor2_1 _11627_ (.A(_05456_),
    .B(_05458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05459_));
 sky130_fd_sc_hd__nor2_1 _11628_ (.A(_05444_),
    .B(_05459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05460_));
 sky130_fd_sc_hd__a21o_1 _11629_ (.A1(_05444_),
    .A2(_05459_),
    .B1(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05461_));
 sky130_fd_sc_hd__nor2_1 _11630_ (.A(_05460_),
    .B(_05461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05462_));
 sky130_fd_sc_hd__buf_2 _11631_ (.A(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05463_));
 sky130_fd_sc_hd__a211o_1 _11632_ (.A1(\sha256cu.data_in_padd[1] ),
    .A2(_05448_),
    .B1(_05462_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05464_));
 sky130_fd_sc_hd__o211a_1 _11633_ (.A1(\sha256cu.iter_processing.w[1] ),
    .A2(_05430_),
    .B1(_05464_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00899_));
 sky130_fd_sc_hd__clkbuf_4 _11634_ (.A(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05465_));
 sky130_fd_sc_hd__or2_1 _11635_ (.A(_05454_),
    .B(_05455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05466_));
 sky130_fd_sc_hd__nand2_1 _11636_ (.A(_05456_),
    .B(_05458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05467_));
 sky130_fd_sc_hd__nand2_1 _11637_ (.A(\sha256cu.msg_scheduler.mreg_9[2] ),
    .B(\sha256cu.msg_scheduler.mreg_0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05468_));
 sky130_fd_sc_hd__or2_1 _11638_ (.A(\sha256cu.msg_scheduler.mreg_9[2] ),
    .B(\sha256cu.msg_scheduler.mreg_0[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05469_));
 sky130_fd_sc_hd__nand2_1 _11639_ (.A(_05468_),
    .B(_05469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05470_));
 sky130_fd_sc_hd__xnor2_1 _11640_ (.A(\sha256cu.msg_scheduler.mreg_1[9] ),
    .B(\sha256cu.msg_scheduler.mreg_1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05471_));
 sky130_fd_sc_hd__xnor2_2 _11641_ (.A(\sha256cu.msg_scheduler.mreg_1[20] ),
    .B(_05471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05472_));
 sky130_fd_sc_hd__xor2_2 _11642_ (.A(_05470_),
    .B(_05472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05473_));
 sky130_fd_sc_hd__a21boi_2 _11643_ (.A1(_05450_),
    .A2(_05453_),
    .B1_N(_05449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05474_));
 sky130_fd_sc_hd__xor2_2 _11644_ (.A(_05473_),
    .B(_05474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05475_));
 sky130_fd_sc_hd__xnor2_1 _11645_ (.A(\sha256cu.msg_scheduler.mreg_14[19] ),
    .B(\sha256cu.msg_scheduler.mreg_14[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05476_));
 sky130_fd_sc_hd__xnor2_1 _11646_ (.A(\sha256cu.msg_scheduler.mreg_14[21] ),
    .B(_05476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05477_));
 sky130_fd_sc_hd__xnor2_1 _11647_ (.A(_05475_),
    .B(_05477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05478_));
 sky130_fd_sc_hd__a21o_1 _11648_ (.A1(_05466_),
    .A2(_05467_),
    .B1(_05478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05479_));
 sky130_fd_sc_hd__nand3_1 _11649_ (.A(_05466_),
    .B(_05467_),
    .C(_05478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05480_));
 sky130_fd_sc_hd__and3_1 _11650_ (.A(_05460_),
    .B(_05479_),
    .C(_05480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05481_));
 sky130_fd_sc_hd__a21oi_1 _11651_ (.A1(_05479_),
    .A2(_05480_),
    .B1(_05460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05482_));
 sky130_fd_sc_hd__nor3_1 _11652_ (.A(_05465_),
    .B(_05481_),
    .C(_05482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05483_));
 sky130_fd_sc_hd__a211o_1 _11653_ (.A1(\sha256cu.data_in_padd[2] ),
    .A2(_05448_),
    .B1(_05483_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05484_));
 sky130_fd_sc_hd__o211a_1 _11654_ (.A1(\sha256cu.iter_processing.w[2] ),
    .A2(_05430_),
    .B1(_05484_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00900_));
 sky130_fd_sc_hd__nand2_1 _11655_ (.A(\sha256cu.msg_scheduler.mreg_9[3] ),
    .B(\sha256cu.msg_scheduler.mreg_0[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05485_));
 sky130_fd_sc_hd__or2_1 _11656_ (.A(\sha256cu.msg_scheduler.mreg_9[3] ),
    .B(\sha256cu.msg_scheduler.mreg_0[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05486_));
 sky130_fd_sc_hd__nand2_1 _11657_ (.A(_05485_),
    .B(_05486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05487_));
 sky130_fd_sc_hd__xnor2_1 _11658_ (.A(\sha256cu.msg_scheduler.mreg_1[10] ),
    .B(\sha256cu.msg_scheduler.mreg_1[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05488_));
 sky130_fd_sc_hd__xnor2_2 _11659_ (.A(\sha256cu.msg_scheduler.mreg_1[21] ),
    .B(_05488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05489_));
 sky130_fd_sc_hd__xor2_1 _11660_ (.A(_05487_),
    .B(_05489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05490_));
 sky130_fd_sc_hd__a21boi_1 _11661_ (.A1(_05469_),
    .A2(_05472_),
    .B1_N(_05468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05491_));
 sky130_fd_sc_hd__or2_1 _11662_ (.A(_05490_),
    .B(_05491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05492_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_05490_),
    .B(_05491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05493_));
 sky130_fd_sc_hd__and2_1 _11664_ (.A(_05492_),
    .B(_05493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05494_));
 sky130_fd_sc_hd__xnor2_1 _11665_ (.A(\sha256cu.msg_scheduler.mreg_14[20] ),
    .B(\sha256cu.msg_scheduler.mreg_14[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05495_));
 sky130_fd_sc_hd__xnor2_1 _11666_ (.A(\sha256cu.msg_scheduler.mreg_14[22] ),
    .B(_05495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05496_));
 sky130_fd_sc_hd__xnor2_1 _11667_ (.A(_05494_),
    .B(_05496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05497_));
 sky130_fd_sc_hd__nor2_1 _11668_ (.A(_05473_),
    .B(_05474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05498_));
 sky130_fd_sc_hd__a21oi_1 _11669_ (.A1(_05475_),
    .A2(_05477_),
    .B1(_05498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05499_));
 sky130_fd_sc_hd__xnor2_1 _11670_ (.A(_05497_),
    .B(_05499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05500_));
 sky130_fd_sc_hd__a21boi_1 _11671_ (.A1(_05460_),
    .A2(_05480_),
    .B1_N(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05501_));
 sky130_fd_sc_hd__or2_1 _11672_ (.A(_05500_),
    .B(_05501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05502_));
 sky130_fd_sc_hd__a21oi_1 _11673_ (.A1(_05500_),
    .A2(_05501_),
    .B1(_05433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05503_));
 sky130_fd_sc_hd__a21o_1 _11674_ (.A1(\sha256cu.data_in_padd[3] ),
    .A2(_05447_),
    .B1(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05504_));
 sky130_fd_sc_hd__a21o_1 _11675_ (.A1(_05502_),
    .A2(_05503_),
    .B1(_05504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05505_));
 sky130_fd_sc_hd__o211a_1 _11676_ (.A1(\sha256cu.iter_processing.w[3] ),
    .A2(_05430_),
    .B1(_05505_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _11677_ (.A(_05497_),
    .B(_05499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05506_));
 sky130_fd_sc_hd__nand2_1 _11678_ (.A(_05494_),
    .B(_05496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05507_));
 sky130_fd_sc_hd__or2_1 _11679_ (.A(\sha256cu.msg_scheduler.mreg_9[4] ),
    .B(\sha256cu.msg_scheduler.mreg_0[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05508_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(\sha256cu.msg_scheduler.mreg_9[4] ),
    .B(\sha256cu.msg_scheduler.mreg_0[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05509_));
 sky130_fd_sc_hd__nand2_1 _11681_ (.A(_05508_),
    .B(_05509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05510_));
 sky130_fd_sc_hd__xnor2_1 _11682_ (.A(\sha256cu.msg_scheduler.mreg_1[11] ),
    .B(\sha256cu.msg_scheduler.mreg_1[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05511_));
 sky130_fd_sc_hd__xnor2_2 _11683_ (.A(\sha256cu.msg_scheduler.mreg_1[22] ),
    .B(_05511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05512_));
 sky130_fd_sc_hd__xor2_1 _11684_ (.A(_05510_),
    .B(_05512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05513_));
 sky130_fd_sc_hd__a21boi_1 _11685_ (.A1(_05486_),
    .A2(_05489_),
    .B1_N(_05485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05514_));
 sky130_fd_sc_hd__or2_1 _11686_ (.A(_05513_),
    .B(_05514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05515_));
 sky130_fd_sc_hd__nand2_1 _11687_ (.A(_05513_),
    .B(_05514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05516_));
 sky130_fd_sc_hd__and2_1 _11688_ (.A(_05515_),
    .B(_05516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05517_));
 sky130_fd_sc_hd__xnor2_1 _11689_ (.A(\sha256cu.msg_scheduler.mreg_14[21] ),
    .B(\sha256cu.msg_scheduler.mreg_14[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05518_));
 sky130_fd_sc_hd__xnor2_1 _11690_ (.A(\sha256cu.msg_scheduler.mreg_14[23] ),
    .B(_05518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05519_));
 sky130_fd_sc_hd__xnor2_1 _11691_ (.A(_05517_),
    .B(_05519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05520_));
 sky130_fd_sc_hd__a21o_1 _11692_ (.A1(_05492_),
    .A2(_05507_),
    .B1(_05520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05521_));
 sky130_fd_sc_hd__nand3_1 _11693_ (.A(_05492_),
    .B(_05507_),
    .C(_05520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_1 _11694_ (.A(_05521_),
    .B(_05522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05523_));
 sky130_fd_sc_hd__a31o_1 _11695_ (.A1(_05506_),
    .A2(_05502_),
    .A3(_05523_),
    .B1(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05524_));
 sky130_fd_sc_hd__a21o_1 _11696_ (.A1(_05506_),
    .A2(_05502_),
    .B1(_05523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05525_));
 sky130_fd_sc_hd__and2b_1 _11697_ (.A_N(_05524_),
    .B(_05525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05526_));
 sky130_fd_sc_hd__a21o_1 _11698_ (.A1(\sha256cu.data_in_padd[4] ),
    .A2(_05448_),
    .B1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05527_));
 sky130_fd_sc_hd__or2_1 _11699_ (.A(\sha256cu.iter_processing.w[4] ),
    .B(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05528_));
 sky130_fd_sc_hd__o211a_1 _11700_ (.A1(_05526_),
    .A2(_05527_),
    .B1(_05528_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00902_));
 sky130_fd_sc_hd__nand2_1 _11701_ (.A(_05517_),
    .B(_05519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05529_));
 sky130_fd_sc_hd__or2_1 _11702_ (.A(\sha256cu.msg_scheduler.mreg_9[5] ),
    .B(\sha256cu.msg_scheduler.mreg_0[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05530_));
 sky130_fd_sc_hd__nand2_1 _11703_ (.A(\sha256cu.msg_scheduler.mreg_9[5] ),
    .B(\sha256cu.msg_scheduler.mreg_0[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_1 _11704_ (.A(_05530_),
    .B(_05531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05532_));
 sky130_fd_sc_hd__xnor2_1 _11705_ (.A(\sha256cu.msg_scheduler.mreg_1[12] ),
    .B(\sha256cu.msg_scheduler.mreg_1[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05533_));
 sky130_fd_sc_hd__xnor2_1 _11706_ (.A(\sha256cu.msg_scheduler.mreg_1[23] ),
    .B(_05533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05534_));
 sky130_fd_sc_hd__xor2_1 _11707_ (.A(_05532_),
    .B(_05534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05535_));
 sky130_fd_sc_hd__a21boi_1 _11708_ (.A1(_05508_),
    .A2(_05512_),
    .B1_N(_05509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05536_));
 sky130_fd_sc_hd__nor2_1 _11709_ (.A(_05535_),
    .B(_05536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05537_));
 sky130_fd_sc_hd__nand2_1 _11710_ (.A(_05535_),
    .B(_05536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05538_));
 sky130_fd_sc_hd__and2b_1 _11711_ (.A_N(_05537_),
    .B(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05539_));
 sky130_fd_sc_hd__xnor2_1 _11712_ (.A(\sha256cu.msg_scheduler.mreg_14[22] ),
    .B(\sha256cu.msg_scheduler.mreg_14[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05540_));
 sky130_fd_sc_hd__xnor2_2 _11713_ (.A(\sha256cu.msg_scheduler.mreg_14[24] ),
    .B(_05540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05541_));
 sky130_fd_sc_hd__xnor2_1 _11714_ (.A(_05539_),
    .B(_05541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05542_));
 sky130_fd_sc_hd__and3_1 _11715_ (.A(_05515_),
    .B(_05529_),
    .C(_05542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05543_));
 sky130_fd_sc_hd__a21o_1 _11716_ (.A1(_05515_),
    .A2(_05529_),
    .B1(_05542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05544_));
 sky130_fd_sc_hd__or2b_1 _11717_ (.A(_05543_),
    .B_N(_05544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05545_));
 sky130_fd_sc_hd__a21oi_1 _11718_ (.A1(_05521_),
    .A2(_05525_),
    .B1(_05545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05546_));
 sky130_fd_sc_hd__a31o_1 _11719_ (.A1(_05521_),
    .A2(_05525_),
    .A3(_05545_),
    .B1(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05547_));
 sky130_fd_sc_hd__nor2_1 _11720_ (.A(_05546_),
    .B(_05547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05548_));
 sky130_fd_sc_hd__a211o_1 _11721_ (.A1(\sha256cu.data_in_padd[5] ),
    .A2(_05448_),
    .B1(_05548_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05549_));
 sky130_fd_sc_hd__o211a_1 _11722_ (.A1(\sha256cu.iter_processing.w[5] ),
    .A2(_05430_),
    .B1(_05549_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00903_));
 sky130_fd_sc_hd__or2_1 _11723_ (.A(\sha256cu.msg_scheduler.mreg_9[6] ),
    .B(\sha256cu.msg_scheduler.mreg_0[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05550_));
 sky130_fd_sc_hd__nand2_1 _11724_ (.A(\sha256cu.msg_scheduler.mreg_9[6] ),
    .B(\sha256cu.msg_scheduler.mreg_0[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_1 _11725_ (.A(_05550_),
    .B(_05551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05552_));
 sky130_fd_sc_hd__xnor2_1 _11726_ (.A(\sha256cu.msg_scheduler.mreg_1[13] ),
    .B(\sha256cu.msg_scheduler.mreg_1[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05553_));
 sky130_fd_sc_hd__xnor2_2 _11727_ (.A(\sha256cu.msg_scheduler.mreg_1[24] ),
    .B(_05553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05554_));
 sky130_fd_sc_hd__xor2_1 _11728_ (.A(_05552_),
    .B(_05554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05555_));
 sky130_fd_sc_hd__a21boi_1 _11729_ (.A1(_05530_),
    .A2(_05534_),
    .B1_N(_05531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05556_));
 sky130_fd_sc_hd__xor2_1 _11730_ (.A(_05555_),
    .B(_05556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05557_));
 sky130_fd_sc_hd__xnor2_1 _11731_ (.A(\sha256cu.msg_scheduler.mreg_14[23] ),
    .B(\sha256cu.msg_scheduler.mreg_14[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05558_));
 sky130_fd_sc_hd__xnor2_1 _11732_ (.A(\sha256cu.msg_scheduler.mreg_14[25] ),
    .B(_05558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_1 _11733_ (.A(_05557_),
    .B(_05559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05560_));
 sky130_fd_sc_hd__or2_1 _11734_ (.A(_05557_),
    .B(_05559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05561_));
 sky130_fd_sc_hd__nand2_1 _11735_ (.A(_05560_),
    .B(_05561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05562_));
 sky130_fd_sc_hd__a21oi_2 _11736_ (.A1(_05538_),
    .A2(_05541_),
    .B1(_05537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05563_));
 sky130_fd_sc_hd__xnor2_1 _11737_ (.A(_05562_),
    .B(_05563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05564_));
 sky130_fd_sc_hd__a21o_1 _11738_ (.A1(_05521_),
    .A2(_05544_),
    .B1(_05543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05565_));
 sky130_fd_sc_hd__o21ai_1 _11739_ (.A1(_05525_),
    .A2(_05545_),
    .B1(_05565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05566_));
 sky130_fd_sc_hd__xor2_1 _11740_ (.A(_05564_),
    .B(_05566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05567_));
 sky130_fd_sc_hd__nor2_1 _11741_ (.A(_05465_),
    .B(_05567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05568_));
 sky130_fd_sc_hd__a211o_1 _11742_ (.A1(\sha256cu.data_in_padd[6] ),
    .A2(_05448_),
    .B1(_05568_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05569_));
 sky130_fd_sc_hd__o211a_1 _11743_ (.A1(\sha256cu.iter_processing.w[6] ),
    .A2(_05430_),
    .B1(_05569_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00904_));
 sky130_fd_sc_hd__or2_1 _11744_ (.A(\sha256cu.msg_scheduler.mreg_9[7] ),
    .B(\sha256cu.msg_scheduler.mreg_0[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05570_));
 sky130_fd_sc_hd__nand2_1 _11745_ (.A(\sha256cu.msg_scheduler.mreg_9[7] ),
    .B(\sha256cu.msg_scheduler.mreg_0[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05571_));
 sky130_fd_sc_hd__nand2_1 _11746_ (.A(_05570_),
    .B(_05571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05572_));
 sky130_fd_sc_hd__xnor2_1 _11747_ (.A(\sha256cu.msg_scheduler.mreg_1[14] ),
    .B(\sha256cu.msg_scheduler.mreg_1[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05573_));
 sky130_fd_sc_hd__xnor2_1 _11748_ (.A(\sha256cu.msg_scheduler.mreg_1[25] ),
    .B(_05573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05574_));
 sky130_fd_sc_hd__xor2_1 _11749_ (.A(_05572_),
    .B(_05574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05575_));
 sky130_fd_sc_hd__a21boi_1 _11750_ (.A1(_05550_),
    .A2(_05554_),
    .B1_N(_05551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05576_));
 sky130_fd_sc_hd__nor2_1 _11751_ (.A(_05575_),
    .B(_05576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05577_));
 sky130_fd_sc_hd__and2_1 _11752_ (.A(_05575_),
    .B(_05576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05578_));
 sky130_fd_sc_hd__nor2_1 _11753_ (.A(_05577_),
    .B(_05578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05579_));
 sky130_fd_sc_hd__xnor2_1 _11754_ (.A(\sha256cu.msg_scheduler.mreg_14[24] ),
    .B(\sha256cu.msg_scheduler.mreg_14[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05580_));
 sky130_fd_sc_hd__xnor2_1 _11755_ (.A(\sha256cu.msg_scheduler.mreg_14[26] ),
    .B(_05580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05581_));
 sky130_fd_sc_hd__xnor2_1 _11756_ (.A(_05579_),
    .B(_05581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05582_));
 sky130_fd_sc_hd__or2_1 _11757_ (.A(_05555_),
    .B(_05556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05583_));
 sky130_fd_sc_hd__nand2_1 _11758_ (.A(_05583_),
    .B(_05560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05584_));
 sky130_fd_sc_hd__xor2_1 _11759_ (.A(_05582_),
    .B(_05584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05585_));
 sky130_fd_sc_hd__nand2_1 _11760_ (.A(_05562_),
    .B(_05563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05586_));
 sky130_fd_sc_hd__nor2_1 _11761_ (.A(_05562_),
    .B(_05563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05587_));
 sky130_fd_sc_hd__a21oi_1 _11762_ (.A1(_05586_),
    .A2(_05566_),
    .B1(_05587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05588_));
 sky130_fd_sc_hd__xnor2_1 _11763_ (.A(_05585_),
    .B(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05589_));
 sky130_fd_sc_hd__nor2_1 _11764_ (.A(_05465_),
    .B(_05589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05590_));
 sky130_fd_sc_hd__a211o_1 _11765_ (.A1(\sha256cu.data_in_padd[7] ),
    .A2(_05448_),
    .B1(_05590_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05591_));
 sky130_fd_sc_hd__o211a_1 _11766_ (.A1(\sha256cu.iter_processing.w[7] ),
    .A2(_05430_),
    .B1(_05591_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00905_));
 sky130_fd_sc_hd__or2_1 _11767_ (.A(_05564_),
    .B(_05585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05592_));
 sky130_fd_sc_hd__or2_1 _11768_ (.A(_05565_),
    .B(_05592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05593_));
 sky130_fd_sc_hd__a2111o_1 _11769_ (.A1(_05506_),
    .A2(_05502_),
    .B1(_05523_),
    .C1(_05545_),
    .D1(_05592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05594_));
 sky130_fd_sc_hd__and2b_1 _11770_ (.A_N(_05582_),
    .B(_05584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05595_));
 sky130_fd_sc_hd__nor2_1 _11771_ (.A(_05587_),
    .B(_05595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05596_));
 sky130_fd_sc_hd__a31o_1 _11772_ (.A1(_05583_),
    .A2(_05560_),
    .A3(_05582_),
    .B1(_05596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05597_));
 sky130_fd_sc_hd__or2_1 _11773_ (.A(\sha256cu.msg_scheduler.mreg_9[8] ),
    .B(\sha256cu.msg_scheduler.mreg_0[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05598_));
 sky130_fd_sc_hd__nand2_1 _11774_ (.A(\sha256cu.msg_scheduler.mreg_9[8] ),
    .B(\sha256cu.msg_scheduler.mreg_0[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05599_));
 sky130_fd_sc_hd__nand2_1 _11775_ (.A(_05598_),
    .B(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05600_));
 sky130_fd_sc_hd__xnor2_1 _11776_ (.A(\sha256cu.msg_scheduler.mreg_1[15] ),
    .B(\sha256cu.msg_scheduler.mreg_1[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05601_));
 sky130_fd_sc_hd__xnor2_1 _11777_ (.A(\sha256cu.msg_scheduler.mreg_1[26] ),
    .B(_05601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05602_));
 sky130_fd_sc_hd__xor2_1 _11778_ (.A(_05600_),
    .B(_05602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05603_));
 sky130_fd_sc_hd__a21boi_1 _11779_ (.A1(_05570_),
    .A2(_05574_),
    .B1_N(_05571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05604_));
 sky130_fd_sc_hd__or2_1 _11780_ (.A(_05603_),
    .B(_05604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05605_));
 sky130_fd_sc_hd__nand2_1 _11781_ (.A(_05603_),
    .B(_05604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05606_));
 sky130_fd_sc_hd__and2_1 _11782_ (.A(_05605_),
    .B(_05606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05607_));
 sky130_fd_sc_hd__xnor2_1 _11783_ (.A(\sha256cu.msg_scheduler.mreg_14[25] ),
    .B(\sha256cu.msg_scheduler.mreg_14[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05608_));
 sky130_fd_sc_hd__xnor2_1 _11784_ (.A(\sha256cu.msg_scheduler.mreg_14[27] ),
    .B(_05608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_1 _11785_ (.A(_05607_),
    .B(_05609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05610_));
 sky130_fd_sc_hd__or2_1 _11786_ (.A(_05607_),
    .B(_05609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05611_));
 sky130_fd_sc_hd__nand2_1 _11787_ (.A(_05610_),
    .B(_05611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05612_));
 sky130_fd_sc_hd__a21oi_1 _11788_ (.A1(_05579_),
    .A2(_05581_),
    .B1(_05577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05613_));
 sky130_fd_sc_hd__xor2_1 _11789_ (.A(_05612_),
    .B(_05613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05614_));
 sky130_fd_sc_hd__inv_2 _11790_ (.A(_05614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05615_));
 sky130_fd_sc_hd__a31o_1 _11791_ (.A1(_05593_),
    .A2(_05594_),
    .A3(_05597_),
    .B1(_05615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05616_));
 sky130_fd_sc_hd__and4_1 _11792_ (.A(_05593_),
    .B(_05594_),
    .C(_05597_),
    .D(_05615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05617_));
 sky130_fd_sc_hd__nor2_1 _11793_ (.A(_05447_),
    .B(_05617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05618_));
 sky130_fd_sc_hd__a221o_1 _11794_ (.A1(\sha256cu.data_in_padd[8] ),
    .A2(_05433_),
    .B1(_05616_),
    .B2(_05618_),
    .C1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05619_));
 sky130_fd_sc_hd__o211a_1 _11795_ (.A1(\sha256cu.iter_processing.w[8] ),
    .A2(_05430_),
    .B1(_05619_),
    .C1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00906_));
 sky130_fd_sc_hd__or2_1 _11796_ (.A(_05612_),
    .B(_05613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05620_));
 sky130_fd_sc_hd__or2_1 _11797_ (.A(\sha256cu.msg_scheduler.mreg_9[9] ),
    .B(\sha256cu.msg_scheduler.mreg_0[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05621_));
 sky130_fd_sc_hd__nand2_1 _11798_ (.A(\sha256cu.msg_scheduler.mreg_9[9] ),
    .B(\sha256cu.msg_scheduler.mreg_0[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05622_));
 sky130_fd_sc_hd__nand2_1 _11799_ (.A(_05621_),
    .B(_05622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05623_));
 sky130_fd_sc_hd__xnor2_1 _11800_ (.A(\sha256cu.msg_scheduler.mreg_1[16] ),
    .B(\sha256cu.msg_scheduler.mreg_1[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05624_));
 sky130_fd_sc_hd__xnor2_1 _11801_ (.A(\sha256cu.msg_scheduler.mreg_1[27] ),
    .B(_05624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05625_));
 sky130_fd_sc_hd__xor2_1 _11802_ (.A(_05623_),
    .B(_05625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05626_));
 sky130_fd_sc_hd__a21boi_1 _11803_ (.A1(_05598_),
    .A2(_05602_),
    .B1_N(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05627_));
 sky130_fd_sc_hd__nor2_1 _11804_ (.A(_05626_),
    .B(_05627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05628_));
 sky130_fd_sc_hd__and2_1 _11805_ (.A(_05626_),
    .B(_05627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05629_));
 sky130_fd_sc_hd__nor2_1 _11806_ (.A(_05628_),
    .B(_05629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05630_));
 sky130_fd_sc_hd__xnor2_1 _11807_ (.A(\sha256cu.msg_scheduler.mreg_14[26] ),
    .B(\sha256cu.msg_scheduler.mreg_14[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05631_));
 sky130_fd_sc_hd__xnor2_1 _11808_ (.A(\sha256cu.msg_scheduler.mreg_14[28] ),
    .B(_05631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05632_));
 sky130_fd_sc_hd__xnor2_1 _11809_ (.A(_05630_),
    .B(_05632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05633_));
 sky130_fd_sc_hd__nand3_1 _11810_ (.A(_05605_),
    .B(_05610_),
    .C(_05633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05634_));
 sky130_fd_sc_hd__a21o_1 _11811_ (.A1(_05605_),
    .A2(_05610_),
    .B1(_05633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05635_));
 sky130_fd_sc_hd__a22o_1 _11812_ (.A1(_05620_),
    .A2(_05616_),
    .B1(_05634_),
    .B2(_05635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05636_));
 sky130_fd_sc_hd__nand4_1 _11813_ (.A(_05620_),
    .B(_05616_),
    .C(_05634_),
    .D(_05635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05637_));
 sky130_fd_sc_hd__a21oi_1 _11814_ (.A1(_05636_),
    .A2(_05637_),
    .B1(_05465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05638_));
 sky130_fd_sc_hd__a211o_1 _11815_ (.A1(\sha256cu.data_in_padd[9] ),
    .A2(_05448_),
    .B1(_05638_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05639_));
 sky130_fd_sc_hd__clkbuf_4 _11816_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05640_));
 sky130_fd_sc_hd__o211a_1 _11817_ (.A1(\sha256cu.iter_processing.w[9] ),
    .A2(_05430_),
    .B1(_05639_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00907_));
 sky130_fd_sc_hd__and2_1 _11818_ (.A(_05620_),
    .B(_05635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05641_));
 sky130_fd_sc_hd__or2_1 _11819_ (.A(\sha256cu.msg_scheduler.mreg_9[10] ),
    .B(\sha256cu.msg_scheduler.mreg_0[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05642_));
 sky130_fd_sc_hd__nand2_1 _11820_ (.A(\sha256cu.msg_scheduler.mreg_9[10] ),
    .B(\sha256cu.msg_scheduler.mreg_0[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05643_));
 sky130_fd_sc_hd__nand2_1 _11821_ (.A(_05642_),
    .B(_05643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05644_));
 sky130_fd_sc_hd__xnor2_1 _11822_ (.A(\sha256cu.msg_scheduler.mreg_1[17] ),
    .B(\sha256cu.msg_scheduler.mreg_1[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05645_));
 sky130_fd_sc_hd__xnor2_1 _11823_ (.A(\sha256cu.msg_scheduler.mreg_1[28] ),
    .B(_05645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05646_));
 sky130_fd_sc_hd__xor2_1 _11824_ (.A(_05644_),
    .B(_05646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05647_));
 sky130_fd_sc_hd__a21boi_1 _11825_ (.A1(_05621_),
    .A2(_05625_),
    .B1_N(_05622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05648_));
 sky130_fd_sc_hd__or2_1 _11826_ (.A(_05647_),
    .B(_05648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05649_));
 sky130_fd_sc_hd__nand2_1 _11827_ (.A(_05647_),
    .B(_05648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05650_));
 sky130_fd_sc_hd__and2_1 _11828_ (.A(_05649_),
    .B(_05650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05651_));
 sky130_fd_sc_hd__xnor2_1 _11829_ (.A(\sha256cu.msg_scheduler.mreg_14[27] ),
    .B(\sha256cu.msg_scheduler.mreg_14[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05652_));
 sky130_fd_sc_hd__xnor2_1 _11830_ (.A(\sha256cu.msg_scheduler.mreg_14[29] ),
    .B(_05652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05653_));
 sky130_fd_sc_hd__nand2_1 _11831_ (.A(_05651_),
    .B(_05653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05654_));
 sky130_fd_sc_hd__or2_1 _11832_ (.A(_05651_),
    .B(_05653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05655_));
 sky130_fd_sc_hd__nand2_1 _11833_ (.A(_05654_),
    .B(_05655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05656_));
 sky130_fd_sc_hd__a21oi_1 _11834_ (.A1(_05630_),
    .A2(_05632_),
    .B1(_05628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05657_));
 sky130_fd_sc_hd__or2_1 _11835_ (.A(_05656_),
    .B(_05657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05658_));
 sky130_fd_sc_hd__nand2_1 _11836_ (.A(_05656_),
    .B(_05657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_1 _11837_ (.A(_05658_),
    .B(_05659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05660_));
 sky130_fd_sc_hd__inv_2 _11838_ (.A(_05634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05661_));
 sky130_fd_sc_hd__a211o_1 _11839_ (.A1(_05616_),
    .A2(_05641_),
    .B1(_05660_),
    .C1(_05661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05662_));
 sky130_fd_sc_hd__a21o_1 _11840_ (.A1(_05616_),
    .A2(_05641_),
    .B1(_05661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05663_));
 sky130_fd_sc_hd__a21oi_1 _11841_ (.A1(_05660_),
    .A2(_05663_),
    .B1(_05465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05664_));
 sky130_fd_sc_hd__a221o_1 _11842_ (.A1(\sha256cu.data_in_padd[10] ),
    .A2(_05433_),
    .B1(_05662_),
    .B2(_05664_),
    .C1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05665_));
 sky130_fd_sc_hd__o211a_1 _11843_ (.A1(\sha256cu.iter_processing.w[10] ),
    .A2(_05430_),
    .B1(_05665_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00908_));
 sky130_fd_sc_hd__clkbuf_4 _11844_ (.A(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05666_));
 sky130_fd_sc_hd__clkbuf_4 _11845_ (.A(_05447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05667_));
 sky130_fd_sc_hd__or2_1 _11846_ (.A(\sha256cu.msg_scheduler.mreg_9[11] ),
    .B(\sha256cu.msg_scheduler.mreg_0[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05668_));
 sky130_fd_sc_hd__nand2_1 _11847_ (.A(\sha256cu.msg_scheduler.mreg_9[11] ),
    .B(\sha256cu.msg_scheduler.mreg_0[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05669_));
 sky130_fd_sc_hd__nand2_1 _11848_ (.A(_05668_),
    .B(_05669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05670_));
 sky130_fd_sc_hd__xnor2_1 _11849_ (.A(\sha256cu.msg_scheduler.mreg_1[18] ),
    .B(\sha256cu.msg_scheduler.mreg_1[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05671_));
 sky130_fd_sc_hd__xnor2_1 _11850_ (.A(\sha256cu.msg_scheduler.mreg_1[29] ),
    .B(_05671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05672_));
 sky130_fd_sc_hd__xor2_1 _11851_ (.A(_05670_),
    .B(_05672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05673_));
 sky130_fd_sc_hd__a21boi_1 _11852_ (.A1(_05642_),
    .A2(_05646_),
    .B1_N(_05643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05674_));
 sky130_fd_sc_hd__nor2_1 _11853_ (.A(_05673_),
    .B(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05675_));
 sky130_fd_sc_hd__and2_1 _11854_ (.A(_05673_),
    .B(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05676_));
 sky130_fd_sc_hd__nor2_1 _11855_ (.A(_05675_),
    .B(_05676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05677_));
 sky130_fd_sc_hd__xnor2_1 _11856_ (.A(\sha256cu.msg_scheduler.mreg_14[28] ),
    .B(\sha256cu.msg_scheduler.mreg_14[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05678_));
 sky130_fd_sc_hd__xnor2_1 _11857_ (.A(\sha256cu.msg_scheduler.mreg_14[30] ),
    .B(_05678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05679_));
 sky130_fd_sc_hd__xnor2_1 _11858_ (.A(_05677_),
    .B(_05679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05680_));
 sky130_fd_sc_hd__and3_1 _11859_ (.A(_05649_),
    .B(_05654_),
    .C(_05680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05681_));
 sky130_fd_sc_hd__a21o_1 _11860_ (.A1(_05649_),
    .A2(_05654_),
    .B1(_05680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05682_));
 sky130_fd_sc_hd__or2b_1 _11861_ (.A(_05681_),
    .B_N(_05682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05683_));
 sky130_fd_sc_hd__a21oi_1 _11862_ (.A1(_05658_),
    .A2(_05662_),
    .B1(_05683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05684_));
 sky130_fd_sc_hd__a31o_1 _11863_ (.A1(_05658_),
    .A2(_05662_),
    .A3(_05683_),
    .B1(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05685_));
 sky130_fd_sc_hd__nor2_1 _11864_ (.A(_05684_),
    .B(_05685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05686_));
 sky130_fd_sc_hd__a211o_1 _11865_ (.A1(\sha256cu.data_in_padd[11] ),
    .A2(_05667_),
    .B1(_05686_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05687_));
 sky130_fd_sc_hd__o211a_1 _11866_ (.A1(\sha256cu.iter_processing.w[11] ),
    .A2(_05666_),
    .B1(_05687_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00909_));
 sky130_fd_sc_hd__or2_1 _11867_ (.A(\sha256cu.msg_scheduler.mreg_9[12] ),
    .B(\sha256cu.msg_scheduler.mreg_0[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05688_));
 sky130_fd_sc_hd__nand2_1 _11868_ (.A(\sha256cu.msg_scheduler.mreg_9[12] ),
    .B(\sha256cu.msg_scheduler.mreg_0[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05689_));
 sky130_fd_sc_hd__nand2_1 _11869_ (.A(_05688_),
    .B(_05689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05690_));
 sky130_fd_sc_hd__xnor2_1 _11870_ (.A(\sha256cu.msg_scheduler.mreg_1[19] ),
    .B(\sha256cu.msg_scheduler.mreg_1[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05691_));
 sky130_fd_sc_hd__xnor2_1 _11871_ (.A(\sha256cu.msg_scheduler.mreg_1[30] ),
    .B(_05691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05692_));
 sky130_fd_sc_hd__xor2_1 _11872_ (.A(_05690_),
    .B(_05692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05693_));
 sky130_fd_sc_hd__a21boi_1 _11873_ (.A1(_05668_),
    .A2(_05672_),
    .B1_N(_05669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05694_));
 sky130_fd_sc_hd__or2_1 _11874_ (.A(_05693_),
    .B(_05694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_1 _11875_ (.A(_05693_),
    .B(_05694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05696_));
 sky130_fd_sc_hd__and2_1 _11876_ (.A(_05695_),
    .B(_05696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05697_));
 sky130_fd_sc_hd__xnor2_1 _11877_ (.A(\sha256cu.msg_scheduler.mreg_14[29] ),
    .B(\sha256cu.msg_scheduler.mreg_14[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05698_));
 sky130_fd_sc_hd__xnor2_1 _11878_ (.A(\sha256cu.msg_scheduler.mreg_14[31] ),
    .B(_05698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05699_));
 sky130_fd_sc_hd__nand2_1 _11879_ (.A(_05697_),
    .B(_05699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05700_));
 sky130_fd_sc_hd__or2_1 _11880_ (.A(_05697_),
    .B(_05699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05701_));
 sky130_fd_sc_hd__nand2_1 _11881_ (.A(_05700_),
    .B(_05701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05702_));
 sky130_fd_sc_hd__a21oi_1 _11882_ (.A1(_05677_),
    .A2(_05679_),
    .B1(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05703_));
 sky130_fd_sc_hd__or2_2 _11883_ (.A(_05702_),
    .B(_05703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05704_));
 sky130_fd_sc_hd__nand2_1 _11884_ (.A(_05702_),
    .B(_05703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05705_));
 sky130_fd_sc_hd__nand2_1 _11885_ (.A(_05704_),
    .B(_05705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05706_));
 sky130_fd_sc_hd__a311o_2 _11886_ (.A1(_05658_),
    .A2(_05662_),
    .A3(_05682_),
    .B1(_05706_),
    .C1(_05681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05707_));
 sky130_fd_sc_hd__a31o_1 _11887_ (.A1(_05658_),
    .A2(_05662_),
    .A3(_05682_),
    .B1(_05681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05708_));
 sky130_fd_sc_hd__a21oi_1 _11888_ (.A1(_05708_),
    .A2(_05706_),
    .B1(_05465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05709_));
 sky130_fd_sc_hd__a221o_1 _11889_ (.A1(\sha256cu.data_in_padd[12] ),
    .A2(_05433_),
    .B1(_05707_),
    .B2(_05709_),
    .C1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05710_));
 sky130_fd_sc_hd__o211a_1 _11890_ (.A1(\sha256cu.iter_processing.w[12] ),
    .A2(_05666_),
    .B1(_05710_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00910_));
 sky130_fd_sc_hd__or2_1 _11891_ (.A(\sha256cu.msg_scheduler.mreg_9[13] ),
    .B(\sha256cu.msg_scheduler.mreg_0[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05711_));
 sky130_fd_sc_hd__nand2_1 _11892_ (.A(\sha256cu.msg_scheduler.mreg_9[13] ),
    .B(\sha256cu.msg_scheduler.mreg_0[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _11893_ (.A(_05711_),
    .B(_05712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05713_));
 sky130_fd_sc_hd__xnor2_1 _11894_ (.A(\sha256cu.msg_scheduler.mreg_1[20] ),
    .B(\sha256cu.msg_scheduler.mreg_1[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05714_));
 sky130_fd_sc_hd__xnor2_1 _11895_ (.A(\sha256cu.msg_scheduler.mreg_1[31] ),
    .B(_05714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05715_));
 sky130_fd_sc_hd__xor2_1 _11896_ (.A(_05713_),
    .B(_05715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05716_));
 sky130_fd_sc_hd__a21boi_1 _11897_ (.A1(_05688_),
    .A2(_05692_),
    .B1_N(_05689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05717_));
 sky130_fd_sc_hd__nor2_1 _11898_ (.A(_05716_),
    .B(_05717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05718_));
 sky130_fd_sc_hd__and2_1 _11899_ (.A(_05716_),
    .B(_05717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05719_));
 sky130_fd_sc_hd__nor2_1 _11900_ (.A(_05718_),
    .B(_05719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05720_));
 sky130_fd_sc_hd__xnor2_1 _11901_ (.A(\sha256cu.msg_scheduler.mreg_14[23] ),
    .B(\sha256cu.msg_scheduler.mreg_14[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05721_));
 sky130_fd_sc_hd__xnor2_1 _11902_ (.A(\sha256cu.msg_scheduler.mreg_14[30] ),
    .B(_05721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05722_));
 sky130_fd_sc_hd__xnor2_1 _11903_ (.A(_05720_),
    .B(_05722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05723_));
 sky130_fd_sc_hd__and3_1 _11904_ (.A(_05695_),
    .B(_05700_),
    .C(_05723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05724_));
 sky130_fd_sc_hd__a21o_1 _11905_ (.A1(_05695_),
    .A2(_05700_),
    .B1(_05723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05725_));
 sky130_fd_sc_hd__or2b_1 _11906_ (.A(_05724_),
    .B_N(_05725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05726_));
 sky130_fd_sc_hd__a21oi_1 _11907_ (.A1(_05704_),
    .A2(_05707_),
    .B1(_05726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05727_));
 sky130_fd_sc_hd__a31o_1 _11908_ (.A1(_05704_),
    .A2(_05707_),
    .A3(_05726_),
    .B1(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05728_));
 sky130_fd_sc_hd__nor2_1 _11909_ (.A(_05727_),
    .B(_05728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05729_));
 sky130_fd_sc_hd__a211o_1 _11910_ (.A1(\sha256cu.data_in_padd[13] ),
    .A2(_05667_),
    .B1(_05729_),
    .C1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05730_));
 sky130_fd_sc_hd__o211a_1 _11911_ (.A1(\sha256cu.iter_processing.w[13] ),
    .A2(_05666_),
    .B1(_05730_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00911_));
 sky130_fd_sc_hd__or2_1 _11912_ (.A(\sha256cu.msg_scheduler.mreg_9[14] ),
    .B(\sha256cu.msg_scheduler.mreg_0[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05731_));
 sky130_fd_sc_hd__nand2_1 _11913_ (.A(\sha256cu.msg_scheduler.mreg_9[14] ),
    .B(\sha256cu.msg_scheduler.mreg_0[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05732_));
 sky130_fd_sc_hd__nand2_1 _11914_ (.A(_05731_),
    .B(_05732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05733_));
 sky130_fd_sc_hd__xnor2_1 _11915_ (.A(\sha256cu.msg_scheduler.mreg_1[17] ),
    .B(\sha256cu.msg_scheduler.mreg_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05734_));
 sky130_fd_sc_hd__xnor2_1 _11916_ (.A(\sha256cu.msg_scheduler.mreg_1[21] ),
    .B(_05734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05735_));
 sky130_fd_sc_hd__xor2_1 _11917_ (.A(_05733_),
    .B(_05735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05736_));
 sky130_fd_sc_hd__a21boi_1 _11918_ (.A1(_05711_),
    .A2(_05715_),
    .B1_N(_05712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05737_));
 sky130_fd_sc_hd__or2_1 _11919_ (.A(_05736_),
    .B(_05737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05738_));
 sky130_fd_sc_hd__nand2_1 _11920_ (.A(_05736_),
    .B(_05737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05739_));
 sky130_fd_sc_hd__and2_1 _11921_ (.A(_05738_),
    .B(_05739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05740_));
 sky130_fd_sc_hd__xnor2_1 _11922_ (.A(\sha256cu.msg_scheduler.mreg_14[24] ),
    .B(\sha256cu.msg_scheduler.mreg_14[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05741_));
 sky130_fd_sc_hd__xnor2_1 _11923_ (.A(\sha256cu.msg_scheduler.mreg_14[31] ),
    .B(_05741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05742_));
 sky130_fd_sc_hd__nand2_1 _11924_ (.A(_05740_),
    .B(_05742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05743_));
 sky130_fd_sc_hd__or2_1 _11925_ (.A(_05740_),
    .B(_05742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05744_));
 sky130_fd_sc_hd__nand2_1 _11926_ (.A(_05743_),
    .B(_05744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05745_));
 sky130_fd_sc_hd__a21oi_1 _11927_ (.A1(_05720_),
    .A2(_05722_),
    .B1(_05718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05746_));
 sky130_fd_sc_hd__or2_2 _11928_ (.A(_05745_),
    .B(_05746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05747_));
 sky130_fd_sc_hd__nand2_1 _11929_ (.A(_05745_),
    .B(_05746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05748_));
 sky130_fd_sc_hd__nand2_1 _11930_ (.A(_05747_),
    .B(_05748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05749_));
 sky130_fd_sc_hd__a311o_4 _11931_ (.A1(_05704_),
    .A2(_05707_),
    .A3(_05725_),
    .B1(_05749_),
    .C1(_05724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05750_));
 sky130_fd_sc_hd__a31o_1 _11932_ (.A1(_05704_),
    .A2(_05707_),
    .A3(_05725_),
    .B1(_05724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05751_));
 sky130_fd_sc_hd__a21oi_1 _11933_ (.A1(_05751_),
    .A2(_05749_),
    .B1(_05433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05752_));
 sky130_fd_sc_hd__a21o_1 _11934_ (.A1(\sha256cu.data_in_padd[14] ),
    .A2(_05447_),
    .B1(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05753_));
 sky130_fd_sc_hd__a21o_1 _11935_ (.A1(_05750_),
    .A2(_05752_),
    .B1(_05753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05754_));
 sky130_fd_sc_hd__o211a_1 _11936_ (.A1(\sha256cu.iter_processing.w[14] ),
    .A2(_05666_),
    .B1(_05754_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00912_));
 sky130_fd_sc_hd__or2_1 _11937_ (.A(\sha256cu.msg_scheduler.mreg_9[15] ),
    .B(\sha256cu.msg_scheduler.mreg_0[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05755_));
 sky130_fd_sc_hd__nand2_1 _11938_ (.A(\sha256cu.msg_scheduler.mreg_9[15] ),
    .B(\sha256cu.msg_scheduler.mreg_0[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05756_));
 sky130_fd_sc_hd__nand2_1 _11939_ (.A(_05755_),
    .B(_05756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05757_));
 sky130_fd_sc_hd__xnor2_1 _11940_ (.A(\sha256cu.msg_scheduler.mreg_1[18] ),
    .B(\sha256cu.msg_scheduler.mreg_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05758_));
 sky130_fd_sc_hd__xnor2_1 _11941_ (.A(\sha256cu.msg_scheduler.mreg_1[22] ),
    .B(_05758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05759_));
 sky130_fd_sc_hd__xor2_1 _11942_ (.A(_05757_),
    .B(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05760_));
 sky130_fd_sc_hd__a21boi_1 _11943_ (.A1(_05731_),
    .A2(_05735_),
    .B1_N(_05732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05761_));
 sky130_fd_sc_hd__nor2_1 _11944_ (.A(_05760_),
    .B(_05761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05762_));
 sky130_fd_sc_hd__and2_1 _11945_ (.A(_05760_),
    .B(_05761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05763_));
 sky130_fd_sc_hd__nor2_1 _11946_ (.A(_05762_),
    .B(_05763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05764_));
 sky130_fd_sc_hd__xnor2_1 _11947_ (.A(\sha256cu.msg_scheduler.mreg_14[2] ),
    .B(\sha256cu.msg_scheduler.mreg_14[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05765_));
 sky130_fd_sc_hd__xnor2_1 _11948_ (.A(\sha256cu.msg_scheduler.mreg_14[25] ),
    .B(_05765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05766_));
 sky130_fd_sc_hd__xnor2_1 _11949_ (.A(_05764_),
    .B(_05766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05767_));
 sky130_fd_sc_hd__and3_1 _11950_ (.A(_05738_),
    .B(_05743_),
    .C(_05767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05768_));
 sky130_fd_sc_hd__a21o_1 _11951_ (.A1(_05738_),
    .A2(_05743_),
    .B1(_05767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05769_));
 sky130_fd_sc_hd__or2b_1 _11952_ (.A(_05768_),
    .B_N(_05769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05770_));
 sky130_fd_sc_hd__a21oi_1 _11953_ (.A1(_05747_),
    .A2(_05750_),
    .B1(_05770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05771_));
 sky130_fd_sc_hd__a31o_1 _11954_ (.A1(_05747_),
    .A2(_05750_),
    .A3(_05770_),
    .B1(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05772_));
 sky130_fd_sc_hd__nor2_1 _11955_ (.A(_05771_),
    .B(_05772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05773_));
 sky130_fd_sc_hd__a211o_1 _11956_ (.A1(\sha256cu.data_in_padd[15] ),
    .A2(_05667_),
    .B1(_05773_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05774_));
 sky130_fd_sc_hd__o211a_1 _11957_ (.A1(\sha256cu.iter_processing.w[15] ),
    .A2(_05666_),
    .B1(_05774_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00913_));
 sky130_fd_sc_hd__a31oi_4 _11958_ (.A1(_05747_),
    .A2(_05750_),
    .A3(_05769_),
    .B1(_05768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05775_));
 sky130_fd_sc_hd__or2_1 _11959_ (.A(\sha256cu.msg_scheduler.mreg_9[16] ),
    .B(\sha256cu.msg_scheduler.mreg_0[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05776_));
 sky130_fd_sc_hd__nand2_1 _11960_ (.A(\sha256cu.msg_scheduler.mreg_9[16] ),
    .B(\sha256cu.msg_scheduler.mreg_0[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_1 _11961_ (.A(_05776_),
    .B(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05778_));
 sky130_fd_sc_hd__xnor2_1 _11962_ (.A(\sha256cu.msg_scheduler.mreg_1[19] ),
    .B(\sha256cu.msg_scheduler.mreg_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05779_));
 sky130_fd_sc_hd__xnor2_1 _11963_ (.A(\sha256cu.msg_scheduler.mreg_1[23] ),
    .B(_05779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05780_));
 sky130_fd_sc_hd__xor2_1 _11964_ (.A(_05778_),
    .B(_05780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05781_));
 sky130_fd_sc_hd__a21boi_2 _11965_ (.A1(_05755_),
    .A2(_05759_),
    .B1_N(_05756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05782_));
 sky130_fd_sc_hd__or2_1 _11966_ (.A(_05781_),
    .B(_05782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05783_));
 sky130_fd_sc_hd__nand2_1 _11967_ (.A(_05781_),
    .B(_05782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05784_));
 sky130_fd_sc_hd__and2_1 _11968_ (.A(_05783_),
    .B(_05784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05785_));
 sky130_fd_sc_hd__xnor2_1 _11969_ (.A(\sha256cu.msg_scheduler.mreg_14[3] ),
    .B(\sha256cu.msg_scheduler.mreg_14[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05786_));
 sky130_fd_sc_hd__xnor2_1 _11970_ (.A(\sha256cu.msg_scheduler.mreg_14[26] ),
    .B(_05786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05787_));
 sky130_fd_sc_hd__nand2_1 _11971_ (.A(_05785_),
    .B(_05787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05788_));
 sky130_fd_sc_hd__or2_1 _11972_ (.A(_05785_),
    .B(_05787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _11973_ (.A(_05788_),
    .B(_05789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05790_));
 sky130_fd_sc_hd__a21oi_1 _11974_ (.A1(_05764_),
    .A2(_05766_),
    .B1(_05762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05791_));
 sky130_fd_sc_hd__or2_1 _11975_ (.A(_05790_),
    .B(_05791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05792_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_05790_),
    .B(_05791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05793_));
 sky130_fd_sc_hd__and2_1 _11977_ (.A(_05792_),
    .B(_05793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05794_));
 sky130_fd_sc_hd__nand2_1 _11978_ (.A(_05775_),
    .B(_05794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05795_));
 sky130_fd_sc_hd__o21a_1 _11979_ (.A1(_05775_),
    .A2(_05794_),
    .B1(_05442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05796_));
 sky130_fd_sc_hd__a221o_1 _11980_ (.A1(\sha256cu.data_in_padd[16] ),
    .A2(_05433_),
    .B1(_05795_),
    .B2(_05796_),
    .C1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05797_));
 sky130_fd_sc_hd__o211a_1 _11981_ (.A1(\sha256cu.iter_processing.w[16] ),
    .A2(_05666_),
    .B1(_05797_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00914_));
 sky130_fd_sc_hd__or2_1 _11982_ (.A(\sha256cu.msg_scheduler.mreg_9[17] ),
    .B(\sha256cu.msg_scheduler.mreg_0[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05798_));
 sky130_fd_sc_hd__nand2_1 _11983_ (.A(\sha256cu.msg_scheduler.mreg_9[17] ),
    .B(\sha256cu.msg_scheduler.mreg_0[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05799_));
 sky130_fd_sc_hd__nand2_1 _11984_ (.A(_05798_),
    .B(_05799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05800_));
 sky130_fd_sc_hd__xnor2_1 _11985_ (.A(\sha256cu.msg_scheduler.mreg_1[20] ),
    .B(\sha256cu.msg_scheduler.mreg_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05801_));
 sky130_fd_sc_hd__xnor2_1 _11986_ (.A(\sha256cu.msg_scheduler.mreg_1[24] ),
    .B(_05801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05802_));
 sky130_fd_sc_hd__xor2_1 _11987_ (.A(_05800_),
    .B(_05802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05803_));
 sky130_fd_sc_hd__a21boi_1 _11988_ (.A1(_05776_),
    .A2(_05780_),
    .B1_N(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05804_));
 sky130_fd_sc_hd__nor2_1 _11989_ (.A(_05803_),
    .B(_05804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05805_));
 sky130_fd_sc_hd__and2_1 _11990_ (.A(_05803_),
    .B(_05804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05806_));
 sky130_fd_sc_hd__nor2_1 _11991_ (.A(_05805_),
    .B(_05806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05807_));
 sky130_fd_sc_hd__xnor2_1 _11992_ (.A(\sha256cu.msg_scheduler.mreg_14[4] ),
    .B(\sha256cu.msg_scheduler.mreg_14[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05808_));
 sky130_fd_sc_hd__xnor2_1 _11993_ (.A(\sha256cu.msg_scheduler.mreg_14[27] ),
    .B(_05808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05809_));
 sky130_fd_sc_hd__xnor2_1 _11994_ (.A(_05807_),
    .B(_05809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05810_));
 sky130_fd_sc_hd__and3_1 _11995_ (.A(_05783_),
    .B(_05788_),
    .C(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05811_));
 sky130_fd_sc_hd__a21o_1 _11996_ (.A1(_05783_),
    .A2(_05788_),
    .B1(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05812_));
 sky130_fd_sc_hd__and2b_1 _11997_ (.A_N(_05811_),
    .B(_05812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05813_));
 sky130_fd_sc_hd__a21oi_1 _11998_ (.A1(_05792_),
    .A2(_05795_),
    .B1(_05813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05814_));
 sky130_fd_sc_hd__and3_1 _11999_ (.A(_05792_),
    .B(_05795_),
    .C(_05813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05815_));
 sky130_fd_sc_hd__o21a_1 _12000_ (.A1(_05814_),
    .A2(_05815_),
    .B1(_05442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05816_));
 sky130_fd_sc_hd__a211o_1 _12001_ (.A1(\sha256cu.data_in_padd[17] ),
    .A2(_05667_),
    .B1(_05816_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05817_));
 sky130_fd_sc_hd__o211a_1 _12002_ (.A1(\sha256cu.iter_processing.w[17] ),
    .A2(_05666_),
    .B1(_05817_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00915_));
 sky130_fd_sc_hd__a21o_1 _12003_ (.A1(_05792_),
    .A2(_05812_),
    .B1(_05811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05818_));
 sky130_fd_sc_hd__and2_1 _12004_ (.A(_05794_),
    .B(_05813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05819_));
 sky130_fd_sc_hd__nand2_1 _12005_ (.A(_05775_),
    .B(_05819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05820_));
 sky130_fd_sc_hd__or2_1 _12006_ (.A(\sha256cu.msg_scheduler.mreg_9[18] ),
    .B(\sha256cu.msg_scheduler.mreg_0[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05821_));
 sky130_fd_sc_hd__nand2_1 _12007_ (.A(\sha256cu.msg_scheduler.mreg_9[18] ),
    .B(\sha256cu.msg_scheduler.mreg_0[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05822_));
 sky130_fd_sc_hd__nand2_1 _12008_ (.A(_05821_),
    .B(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05823_));
 sky130_fd_sc_hd__xnor2_1 _12009_ (.A(\sha256cu.msg_scheduler.mreg_1[21] ),
    .B(\sha256cu.msg_scheduler.mreg_1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05824_));
 sky130_fd_sc_hd__xnor2_1 _12010_ (.A(\sha256cu.msg_scheduler.mreg_1[25] ),
    .B(_05824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05825_));
 sky130_fd_sc_hd__xor2_1 _12011_ (.A(_05823_),
    .B(_05825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05826_));
 sky130_fd_sc_hd__a21boi_1 _12012_ (.A1(_05798_),
    .A2(_05802_),
    .B1_N(_05799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05827_));
 sky130_fd_sc_hd__or2_1 _12013_ (.A(_05826_),
    .B(_05827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05828_));
 sky130_fd_sc_hd__nand2_1 _12014_ (.A(_05826_),
    .B(_05827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05829_));
 sky130_fd_sc_hd__and2_1 _12015_ (.A(_05828_),
    .B(_05829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05830_));
 sky130_fd_sc_hd__xnor2_1 _12016_ (.A(\sha256cu.msg_scheduler.mreg_14[5] ),
    .B(\sha256cu.msg_scheduler.mreg_14[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05831_));
 sky130_fd_sc_hd__xnor2_1 _12017_ (.A(\sha256cu.msg_scheduler.mreg_14[28] ),
    .B(_05831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05832_));
 sky130_fd_sc_hd__nand2_1 _12018_ (.A(_05830_),
    .B(_05832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05833_));
 sky130_fd_sc_hd__or2_1 _12019_ (.A(_05830_),
    .B(_05832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05834_));
 sky130_fd_sc_hd__nand2_1 _12020_ (.A(_05833_),
    .B(_05834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05835_));
 sky130_fd_sc_hd__a21oi_1 _12021_ (.A1(_05807_),
    .A2(_05809_),
    .B1(_05805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05836_));
 sky130_fd_sc_hd__nor2_1 _12022_ (.A(_05835_),
    .B(_05836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05837_));
 sky130_fd_sc_hd__inv_2 _12023_ (.A(_05837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_1 _12024_ (.A(_05835_),
    .B(_05836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05839_));
 sky130_fd_sc_hd__nand2_1 _12025_ (.A(_05838_),
    .B(_05839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05840_));
 sky130_fd_sc_hd__a21o_1 _12026_ (.A1(_05818_),
    .A2(_05820_),
    .B1(_05840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05841_));
 sky130_fd_sc_hd__a31oi_1 _12027_ (.A1(_05840_),
    .A2(_05818_),
    .A3(_05820_),
    .B1(_05433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05842_));
 sky130_fd_sc_hd__a21o_1 _12028_ (.A1(\sha256cu.data_in_padd[18] ),
    .A2(_05447_),
    .B1(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05843_));
 sky130_fd_sc_hd__a21o_1 _12029_ (.A1(_05841_),
    .A2(_05842_),
    .B1(_05843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05844_));
 sky130_fd_sc_hd__o211a_1 _12030_ (.A1(\sha256cu.iter_processing.w[18] ),
    .A2(_05666_),
    .B1(_05844_),
    .C1(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00916_));
 sky130_fd_sc_hd__or2_1 _12031_ (.A(\sha256cu.msg_scheduler.mreg_9[19] ),
    .B(\sha256cu.msg_scheduler.mreg_0[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05845_));
 sky130_fd_sc_hd__nand2_1 _12032_ (.A(\sha256cu.msg_scheduler.mreg_9[19] ),
    .B(\sha256cu.msg_scheduler.mreg_0[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_05845_),
    .B(_05846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05847_));
 sky130_fd_sc_hd__xnor2_1 _12034_ (.A(\sha256cu.msg_scheduler.mreg_1[22] ),
    .B(\sha256cu.msg_scheduler.mreg_1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05848_));
 sky130_fd_sc_hd__xnor2_1 _12035_ (.A(\sha256cu.msg_scheduler.mreg_1[26] ),
    .B(_05848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05849_));
 sky130_fd_sc_hd__xor2_1 _12036_ (.A(_05847_),
    .B(_05849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05850_));
 sky130_fd_sc_hd__a21boi_1 _12037_ (.A1(_05821_),
    .A2(_05825_),
    .B1_N(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05851_));
 sky130_fd_sc_hd__nor2_1 _12038_ (.A(_05850_),
    .B(_05851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05852_));
 sky130_fd_sc_hd__and2_1 _12039_ (.A(_05850_),
    .B(_05851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05853_));
 sky130_fd_sc_hd__nor2_1 _12040_ (.A(_05852_),
    .B(_05853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05854_));
 sky130_fd_sc_hd__xnor2_1 _12041_ (.A(\sha256cu.msg_scheduler.mreg_14[6] ),
    .B(\sha256cu.msg_scheduler.mreg_14[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05855_));
 sky130_fd_sc_hd__xnor2_1 _12042_ (.A(\sha256cu.msg_scheduler.mreg_14[29] ),
    .B(_05855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05856_));
 sky130_fd_sc_hd__xnor2_1 _12043_ (.A(_05854_),
    .B(_05856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05857_));
 sky130_fd_sc_hd__and3_1 _12044_ (.A(_05828_),
    .B(_05833_),
    .C(_05857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05858_));
 sky130_fd_sc_hd__a21o_1 _12045_ (.A1(_05828_),
    .A2(_05833_),
    .B1(_05857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05859_));
 sky130_fd_sc_hd__and2b_1 _12046_ (.A_N(_05858_),
    .B(_05859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05860_));
 sky130_fd_sc_hd__inv_2 _12047_ (.A(_05860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05861_));
 sky130_fd_sc_hd__a21oi_1 _12048_ (.A1(_05838_),
    .A2(_05841_),
    .B1(_05861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05862_));
 sky130_fd_sc_hd__a31o_1 _12049_ (.A1(_05838_),
    .A2(_05841_),
    .A3(_05861_),
    .B1(_05465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05863_));
 sky130_fd_sc_hd__a21oi_1 _12050_ (.A1(\sha256cu.data_in_padd[19] ),
    .A2(_05667_),
    .B1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05864_));
 sky130_fd_sc_hd__o21ai_1 _12051_ (.A1(_05862_),
    .A2(_05863_),
    .B1(_05864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05865_));
 sky130_fd_sc_hd__clkbuf_4 _12052_ (.A(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05866_));
 sky130_fd_sc_hd__o211a_1 _12053_ (.A1(\sha256cu.iter_processing.w[19] ),
    .A2(_05666_),
    .B1(_05865_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00917_));
 sky130_fd_sc_hd__or2_1 _12054_ (.A(\sha256cu.msg_scheduler.mreg_9[20] ),
    .B(\sha256cu.msg_scheduler.mreg_0[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05867_));
 sky130_fd_sc_hd__nand2_1 _12055_ (.A(\sha256cu.msg_scheduler.mreg_9[20] ),
    .B(\sha256cu.msg_scheduler.mreg_0[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05868_));
 sky130_fd_sc_hd__nand2_1 _12056_ (.A(_05867_),
    .B(_05868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05869_));
 sky130_fd_sc_hd__xnor2_1 _12057_ (.A(\sha256cu.msg_scheduler.mreg_1[23] ),
    .B(\sha256cu.msg_scheduler.mreg_1[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05870_));
 sky130_fd_sc_hd__xnor2_1 _12058_ (.A(\sha256cu.msg_scheduler.mreg_1[27] ),
    .B(_05870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05871_));
 sky130_fd_sc_hd__xor2_1 _12059_ (.A(_05869_),
    .B(_05871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05872_));
 sky130_fd_sc_hd__a21boi_1 _12060_ (.A1(_05845_),
    .A2(_05849_),
    .B1_N(_05846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05873_));
 sky130_fd_sc_hd__or2_1 _12061_ (.A(_05872_),
    .B(_05873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05874_));
 sky130_fd_sc_hd__nand2_1 _12062_ (.A(_05872_),
    .B(_05873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05875_));
 sky130_fd_sc_hd__and2_1 _12063_ (.A(_05874_),
    .B(_05875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05876_));
 sky130_fd_sc_hd__xnor2_1 _12064_ (.A(\sha256cu.msg_scheduler.mreg_14[7] ),
    .B(\sha256cu.msg_scheduler.mreg_14[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05877_));
 sky130_fd_sc_hd__xnor2_1 _12065_ (.A(\sha256cu.msg_scheduler.mreg_14[30] ),
    .B(_05877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_1 _12066_ (.A(_05876_),
    .B(_05878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05879_));
 sky130_fd_sc_hd__or2_1 _12067_ (.A(_05876_),
    .B(_05878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05880_));
 sky130_fd_sc_hd__nand2_1 _12068_ (.A(_05879_),
    .B(_05880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05881_));
 sky130_fd_sc_hd__a21oi_1 _12069_ (.A1(_05854_),
    .A2(_05856_),
    .B1(_05852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05882_));
 sky130_fd_sc_hd__or2_1 _12070_ (.A(_05881_),
    .B(_05882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05883_));
 sky130_fd_sc_hd__nand2_1 _12071_ (.A(_05881_),
    .B(_05882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05884_));
 sky130_fd_sc_hd__and2_1 _12072_ (.A(_05883_),
    .B(_05884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05885_));
 sky130_fd_sc_hd__nand3b_1 _12073_ (.A_N(_05840_),
    .B(_05819_),
    .C(_05860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05886_));
 sky130_fd_sc_hd__inv_2 _12074_ (.A(_05886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05887_));
 sky130_fd_sc_hd__o32a_1 _12075_ (.A1(_05840_),
    .A2(_05818_),
    .A3(_05861_),
    .B1(_05858_),
    .B2(_05838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05888_));
 sky130_fd_sc_hd__and2_1 _12076_ (.A(_05859_),
    .B(_05888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05889_));
 sky130_fd_sc_hd__a21bo_1 _12077_ (.A1(_05775_),
    .A2(_05887_),
    .B1_N(_05889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05890_));
 sky130_fd_sc_hd__nand2_1 _12078_ (.A(_05885_),
    .B(_05890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05891_));
 sky130_fd_sc_hd__o211a_1 _12079_ (.A1(_05885_),
    .A2(_05890_),
    .B1(_05891_),
    .C1(_05442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05892_));
 sky130_fd_sc_hd__a211o_1 _12080_ (.A1(\sha256cu.data_in_padd[20] ),
    .A2(_05667_),
    .B1(_05892_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05893_));
 sky130_fd_sc_hd__o211a_1 _12081_ (.A1(\sha256cu.iter_processing.w[20] ),
    .A2(_05666_),
    .B1(_05893_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00918_));
 sky130_fd_sc_hd__clkbuf_4 _12082_ (.A(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05894_));
 sky130_fd_sc_hd__or2_1 _12083_ (.A(\sha256cu.msg_scheduler.mreg_9[21] ),
    .B(\sha256cu.msg_scheduler.mreg_0[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05895_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(\sha256cu.msg_scheduler.mreg_9[21] ),
    .B(\sha256cu.msg_scheduler.mreg_0[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05896_));
 sky130_fd_sc_hd__nand2_1 _12085_ (.A(_05895_),
    .B(_05896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05897_));
 sky130_fd_sc_hd__xnor2_1 _12086_ (.A(\sha256cu.msg_scheduler.mreg_1[24] ),
    .B(\sha256cu.msg_scheduler.mreg_1[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05898_));
 sky130_fd_sc_hd__xnor2_1 _12087_ (.A(\sha256cu.msg_scheduler.mreg_1[28] ),
    .B(_05898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05899_));
 sky130_fd_sc_hd__xor2_1 _12088_ (.A(_05897_),
    .B(_05899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05900_));
 sky130_fd_sc_hd__a21boi_1 _12089_ (.A1(_05867_),
    .A2(_05871_),
    .B1_N(_05868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05901_));
 sky130_fd_sc_hd__nor2_1 _12090_ (.A(_05900_),
    .B(_05901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05902_));
 sky130_fd_sc_hd__and2_1 _12091_ (.A(_05900_),
    .B(_05901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05903_));
 sky130_fd_sc_hd__nor2_1 _12092_ (.A(_05902_),
    .B(_05903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05904_));
 sky130_fd_sc_hd__xnor2_1 _12093_ (.A(\sha256cu.msg_scheduler.mreg_14[8] ),
    .B(\sha256cu.msg_scheduler.mreg_14[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05905_));
 sky130_fd_sc_hd__xnor2_1 _12094_ (.A(\sha256cu.msg_scheduler.mreg_14[31] ),
    .B(_05905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05906_));
 sky130_fd_sc_hd__xnor2_1 _12095_ (.A(_05904_),
    .B(_05906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05907_));
 sky130_fd_sc_hd__and3_1 _12096_ (.A(_05874_),
    .B(_05879_),
    .C(_05907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05908_));
 sky130_fd_sc_hd__a21o_1 _12097_ (.A1(_05874_),
    .A2(_05879_),
    .B1(_05907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05909_));
 sky130_fd_sc_hd__and2b_1 _12098_ (.A_N(_05908_),
    .B(_05909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05910_));
 sky130_fd_sc_hd__a21oi_1 _12099_ (.A1(_05883_),
    .A2(_05891_),
    .B1(_05910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05911_));
 sky130_fd_sc_hd__and3_1 _12100_ (.A(_05883_),
    .B(_05891_),
    .C(_05910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05912_));
 sky130_fd_sc_hd__or2_1 _12101_ (.A(_05911_),
    .B(_05912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05913_));
 sky130_fd_sc_hd__a21o_1 _12102_ (.A1(\sha256cu.data_in_padd[21] ),
    .A2(_05447_),
    .B1(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05914_));
 sky130_fd_sc_hd__a21o_1 _12103_ (.A1(_05442_),
    .A2(_05913_),
    .B1(_05914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05915_));
 sky130_fd_sc_hd__o211a_1 _12104_ (.A1(\sha256cu.iter_processing.w[21] ),
    .A2(_05894_),
    .B1(_05915_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00919_));
 sky130_fd_sc_hd__or2_1 _12105_ (.A(\sha256cu.msg_scheduler.mreg_9[22] ),
    .B(\sha256cu.msg_scheduler.mreg_0[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05916_));
 sky130_fd_sc_hd__nand2_1 _12106_ (.A(\sha256cu.msg_scheduler.mreg_9[22] ),
    .B(\sha256cu.msg_scheduler.mreg_0[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05917_));
 sky130_fd_sc_hd__nand2_1 _12107_ (.A(_05916_),
    .B(_05917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05918_));
 sky130_fd_sc_hd__xnor2_1 _12108_ (.A(\sha256cu.msg_scheduler.mreg_1[25] ),
    .B(\sha256cu.msg_scheduler.mreg_1[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05919_));
 sky130_fd_sc_hd__xnor2_1 _12109_ (.A(\sha256cu.msg_scheduler.mreg_1[29] ),
    .B(_05919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05920_));
 sky130_fd_sc_hd__xor2_1 _12110_ (.A(_05918_),
    .B(_05920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05921_));
 sky130_fd_sc_hd__a21boi_1 _12111_ (.A1(_05895_),
    .A2(_05899_),
    .B1_N(_05896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05922_));
 sky130_fd_sc_hd__or2_1 _12112_ (.A(_05921_),
    .B(_05922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05923_));
 sky130_fd_sc_hd__nand2_1 _12113_ (.A(_05921_),
    .B(_05922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05924_));
 sky130_fd_sc_hd__and2_1 _12114_ (.A(_05923_),
    .B(_05924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05925_));
 sky130_fd_sc_hd__xor2_1 _12115_ (.A(\sha256cu.msg_scheduler.mreg_14[9] ),
    .B(\sha256cu.msg_scheduler.mreg_14[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05926_));
 sky130_fd_sc_hd__nand2_1 _12116_ (.A(_05925_),
    .B(_05926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05927_));
 sky130_fd_sc_hd__or2_1 _12117_ (.A(_05925_),
    .B(_05926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05928_));
 sky130_fd_sc_hd__nand2_1 _12118_ (.A(_05927_),
    .B(_05928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05929_));
 sky130_fd_sc_hd__a21oi_1 _12119_ (.A1(_05904_),
    .A2(_05906_),
    .B1(_05902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05930_));
 sky130_fd_sc_hd__nor2_1 _12120_ (.A(_05929_),
    .B(_05930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05931_));
 sky130_fd_sc_hd__and2_1 _12121_ (.A(_05929_),
    .B(_05930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05932_));
 sky130_fd_sc_hd__or2_1 _12122_ (.A(_05931_),
    .B(_05932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05933_));
 sky130_fd_sc_hd__inv_2 _12123_ (.A(_05933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05934_));
 sky130_fd_sc_hd__and2_1 _12124_ (.A(_05885_),
    .B(_05910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05935_));
 sky130_fd_sc_hd__a21o_1 _12125_ (.A1(_05883_),
    .A2(_05909_),
    .B1(_05908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05936_));
 sky130_fd_sc_hd__a21bo_1 _12126_ (.A1(_05890_),
    .A2(_05935_),
    .B1_N(_05936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05937_));
 sky130_fd_sc_hd__xnor2_1 _12127_ (.A(_05934_),
    .B(_05937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05938_));
 sky130_fd_sc_hd__nor2_1 _12128_ (.A(_05465_),
    .B(_05938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05939_));
 sky130_fd_sc_hd__a211o_1 _12129_ (.A1(\sha256cu.data_in_padd[22] ),
    .A2(_05667_),
    .B1(_05939_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05940_));
 sky130_fd_sc_hd__o211a_1 _12130_ (.A1(\sha256cu.iter_processing.w[22] ),
    .A2(_05894_),
    .B1(_05940_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00920_));
 sky130_fd_sc_hd__or2_1 _12131_ (.A(\sha256cu.msg_scheduler.mreg_9[23] ),
    .B(\sha256cu.msg_scheduler.mreg_0[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05941_));
 sky130_fd_sc_hd__nand2_1 _12132_ (.A(\sha256cu.msg_scheduler.mreg_9[23] ),
    .B(\sha256cu.msg_scheduler.mreg_0[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05942_));
 sky130_fd_sc_hd__nand2_1 _12133_ (.A(_05941_),
    .B(_05942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05943_));
 sky130_fd_sc_hd__xnor2_1 _12134_ (.A(\sha256cu.msg_scheduler.mreg_1[26] ),
    .B(\sha256cu.msg_scheduler.mreg_1[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05944_));
 sky130_fd_sc_hd__xnor2_1 _12135_ (.A(\sha256cu.msg_scheduler.mreg_1[30] ),
    .B(_05944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05945_));
 sky130_fd_sc_hd__xor2_1 _12136_ (.A(_05943_),
    .B(_05945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05946_));
 sky130_fd_sc_hd__a21boi_1 _12137_ (.A1(_05916_),
    .A2(_05920_),
    .B1_N(_05917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05947_));
 sky130_fd_sc_hd__nor2_1 _12138_ (.A(_05946_),
    .B(_05947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05948_));
 sky130_fd_sc_hd__and2_1 _12139_ (.A(_05946_),
    .B(_05947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05949_));
 sky130_fd_sc_hd__nor2_1 _12140_ (.A(_05948_),
    .B(_05949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05950_));
 sky130_fd_sc_hd__xor2_1 _12141_ (.A(\sha256cu.msg_scheduler.mreg_14[10] ),
    .B(\sha256cu.msg_scheduler.mreg_14[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05951_));
 sky130_fd_sc_hd__xnor2_1 _12142_ (.A(_05950_),
    .B(_05951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05952_));
 sky130_fd_sc_hd__nand3_1 _12143_ (.A(_05923_),
    .B(_05927_),
    .C(_05952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05953_));
 sky130_fd_sc_hd__inv_2 _12144_ (.A(_05953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05954_));
 sky130_fd_sc_hd__a21oi_1 _12145_ (.A1(_05923_),
    .A2(_05927_),
    .B1(_05952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05955_));
 sky130_fd_sc_hd__nor2_1 _12146_ (.A(_05954_),
    .B(_05955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05956_));
 sky130_fd_sc_hd__a21oi_1 _12147_ (.A1(_05934_),
    .A2(_05937_),
    .B1(_05931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05957_));
 sky130_fd_sc_hd__xnor2_1 _12148_ (.A(_05956_),
    .B(_05957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05958_));
 sky130_fd_sc_hd__a21o_1 _12149_ (.A1(\sha256cu.data_in_padd[23] ),
    .A2(_05447_),
    .B1(_04692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05959_));
 sky130_fd_sc_hd__a21o_1 _12150_ (.A1(_05442_),
    .A2(_05958_),
    .B1(_05959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05960_));
 sky130_fd_sc_hd__o211a_1 _12151_ (.A1(\sha256cu.iter_processing.w[23] ),
    .A2(_05894_),
    .B1(_05960_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00921_));
 sky130_fd_sc_hd__nand3_1 _12152_ (.A(_05934_),
    .B(_05935_),
    .C(_05956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05961_));
 sky130_fd_sc_hd__or2_1 _12153_ (.A(_05886_),
    .B(_05961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05962_));
 sky130_fd_sc_hd__a311o_1 _12154_ (.A1(_05747_),
    .A2(_05750_),
    .A3(_05769_),
    .B1(_05962_),
    .C1(_05768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05963_));
 sky130_fd_sc_hd__or3b_1 _12155_ (.A(_05933_),
    .B(_05936_),
    .C_N(_05956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05964_));
 sky130_fd_sc_hd__a21oi_1 _12156_ (.A1(_05931_),
    .A2(_05953_),
    .B1(_05955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05965_));
 sky130_fd_sc_hd__o211a_1 _12157_ (.A1(_05889_),
    .A2(_05961_),
    .B1(_05964_),
    .C1(_05965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05966_));
 sky130_fd_sc_hd__and2_1 _12158_ (.A(_05963_),
    .B(_05966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05967_));
 sky130_fd_sc_hd__or2_1 _12159_ (.A(\sha256cu.msg_scheduler.mreg_9[24] ),
    .B(\sha256cu.msg_scheduler.mreg_0[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05968_));
 sky130_fd_sc_hd__nand2_1 _12160_ (.A(\sha256cu.msg_scheduler.mreg_9[24] ),
    .B(\sha256cu.msg_scheduler.mreg_0[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2_1 _12161_ (.A(_05968_),
    .B(_05969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05970_));
 sky130_fd_sc_hd__xnor2_1 _12162_ (.A(\sha256cu.msg_scheduler.mreg_1[27] ),
    .B(\sha256cu.msg_scheduler.mreg_1[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05971_));
 sky130_fd_sc_hd__xnor2_1 _12163_ (.A(\sha256cu.msg_scheduler.mreg_1[31] ),
    .B(_05971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05972_));
 sky130_fd_sc_hd__xor2_1 _12164_ (.A(_05970_),
    .B(_05972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05973_));
 sky130_fd_sc_hd__a21boi_1 _12165_ (.A1(_05941_),
    .A2(_05945_),
    .B1_N(_05942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05974_));
 sky130_fd_sc_hd__or2_1 _12166_ (.A(_05973_),
    .B(_05974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05975_));
 sky130_fd_sc_hd__nand2_1 _12167_ (.A(_05973_),
    .B(_05974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05976_));
 sky130_fd_sc_hd__nand2_1 _12168_ (.A(_05975_),
    .B(_05976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05977_));
 sky130_fd_sc_hd__xor2_1 _12169_ (.A(\sha256cu.msg_scheduler.mreg_14[11] ),
    .B(\sha256cu.msg_scheduler.mreg_14[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05978_));
 sky130_fd_sc_hd__xor2_1 _12170_ (.A(_05977_),
    .B(_05978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05979_));
 sky130_fd_sc_hd__a21oi_1 _12171_ (.A1(_05950_),
    .A2(_05951_),
    .B1(_05948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05980_));
 sky130_fd_sc_hd__or2_1 _12172_ (.A(_05979_),
    .B(_05980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05981_));
 sky130_fd_sc_hd__nand2_1 _12173_ (.A(_05979_),
    .B(_05980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05982_));
 sky130_fd_sc_hd__and2_1 _12174_ (.A(_05981_),
    .B(_05982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05983_));
 sky130_fd_sc_hd__inv_2 _12175_ (.A(_05983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05984_));
 sky130_fd_sc_hd__a21oi_1 _12176_ (.A1(_05967_),
    .A2(_05984_),
    .B1(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05985_));
 sky130_fd_sc_hd__o21a_1 _12177_ (.A1(_05967_),
    .A2(_05984_),
    .B1(_05985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05986_));
 sky130_fd_sc_hd__a211o_1 _12178_ (.A1(\sha256cu.data_in_padd[24] ),
    .A2(_05667_),
    .B1(_05986_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05987_));
 sky130_fd_sc_hd__o211a_1 _12179_ (.A1(\sha256cu.iter_processing.w[24] ),
    .A2(_05894_),
    .B1(_05987_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00922_));
 sky130_fd_sc_hd__or2b_1 _12180_ (.A(_05977_),
    .B_N(_05978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05988_));
 sky130_fd_sc_hd__or2_1 _12181_ (.A(\sha256cu.msg_scheduler.mreg_9[25] ),
    .B(\sha256cu.msg_scheduler.mreg_0[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05989_));
 sky130_fd_sc_hd__nand2_1 _12182_ (.A(\sha256cu.msg_scheduler.mreg_9[25] ),
    .B(\sha256cu.msg_scheduler.mreg_0[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2_1 _12183_ (.A(_05989_),
    .B(_05990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05991_));
 sky130_fd_sc_hd__xnor2_1 _12184_ (.A(\sha256cu.msg_scheduler.mreg_1[11] ),
    .B(\sha256cu.msg_scheduler.mreg_1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05992_));
 sky130_fd_sc_hd__xnor2_1 _12185_ (.A(\sha256cu.msg_scheduler.mreg_1[28] ),
    .B(_05992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05993_));
 sky130_fd_sc_hd__xor2_1 _12186_ (.A(_05991_),
    .B(_05993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05994_));
 sky130_fd_sc_hd__a21boi_1 _12187_ (.A1(_05968_),
    .A2(_05972_),
    .B1_N(_05969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05995_));
 sky130_fd_sc_hd__or2_1 _12188_ (.A(_05994_),
    .B(_05995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05996_));
 sky130_fd_sc_hd__nand2_1 _12189_ (.A(_05994_),
    .B(_05995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05997_));
 sky130_fd_sc_hd__and2_1 _12190_ (.A(_05996_),
    .B(_05997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05998_));
 sky130_fd_sc_hd__xor2_1 _12191_ (.A(\sha256cu.msg_scheduler.mreg_14[12] ),
    .B(\sha256cu.msg_scheduler.mreg_14[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05999_));
 sky130_fd_sc_hd__nand2_1 _12192_ (.A(_05998_),
    .B(_05999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06000_));
 sky130_fd_sc_hd__or2_1 _12193_ (.A(_05998_),
    .B(_05999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06001_));
 sky130_fd_sc_hd__nand2_1 _12194_ (.A(_06000_),
    .B(_06001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06002_));
 sky130_fd_sc_hd__and3_1 _12195_ (.A(_05975_),
    .B(_05988_),
    .C(_06002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06003_));
 sky130_fd_sc_hd__a21o_1 _12196_ (.A1(_05975_),
    .A2(_05988_),
    .B1(_06002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06004_));
 sky130_fd_sc_hd__and2b_1 _12197_ (.A_N(_06003_),
    .B(_06004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06005_));
 sky130_fd_sc_hd__o21ai_1 _12198_ (.A1(_05967_),
    .A2(_05984_),
    .B1(_05981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2_1 _12199_ (.A(_06005_),
    .B(_06006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06007_));
 sky130_fd_sc_hd__o211a_1 _12200_ (.A1(_06005_),
    .A2(_06006_),
    .B1(_06007_),
    .C1(_05442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06008_));
 sky130_fd_sc_hd__a211o_1 _12201_ (.A1(\sha256cu.data_in_padd[25] ),
    .A2(_05667_),
    .B1(_06008_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06009_));
 sky130_fd_sc_hd__o211a_1 _12202_ (.A1(\sha256cu.iter_processing.w[25] ),
    .A2(_05894_),
    .B1(_06009_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00923_));
 sky130_fd_sc_hd__or2_1 _12203_ (.A(\sha256cu.msg_scheduler.mreg_9[26] ),
    .B(\sha256cu.msg_scheduler.mreg_0[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06010_));
 sky130_fd_sc_hd__nand2_1 _12204_ (.A(\sha256cu.msg_scheduler.mreg_9[26] ),
    .B(\sha256cu.msg_scheduler.mreg_0[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(_06010_),
    .B(_06011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06012_));
 sky130_fd_sc_hd__xnor2_1 _12206_ (.A(\sha256cu.msg_scheduler.mreg_1[12] ),
    .B(\sha256cu.msg_scheduler.mreg_1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06013_));
 sky130_fd_sc_hd__xnor2_1 _12207_ (.A(\sha256cu.msg_scheduler.mreg_1[29] ),
    .B(_06013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06014_));
 sky130_fd_sc_hd__xor2_1 _12208_ (.A(_06012_),
    .B(_06014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06015_));
 sky130_fd_sc_hd__a21boi_1 _12209_ (.A1(_05989_),
    .A2(_05993_),
    .B1_N(_05990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06016_));
 sky130_fd_sc_hd__or2_1 _12210_ (.A(_06015_),
    .B(_06016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06017_));
 sky130_fd_sc_hd__nand2_1 _12211_ (.A(_06015_),
    .B(_06016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06018_));
 sky130_fd_sc_hd__and2_1 _12212_ (.A(_06017_),
    .B(_06018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06019_));
 sky130_fd_sc_hd__xor2_1 _12213_ (.A(\sha256cu.msg_scheduler.mreg_14[13] ),
    .B(\sha256cu.msg_scheduler.mreg_14[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06020_));
 sky130_fd_sc_hd__nand2_1 _12214_ (.A(_06019_),
    .B(_06020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06021_));
 sky130_fd_sc_hd__or2_1 _12215_ (.A(_06019_),
    .B(_06020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06022_));
 sky130_fd_sc_hd__nand2_1 _12216_ (.A(_06021_),
    .B(_06022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06023_));
 sky130_fd_sc_hd__a21oi_2 _12217_ (.A1(_05996_),
    .A2(_06000_),
    .B1(_06023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06024_));
 sky130_fd_sc_hd__and3_1 _12218_ (.A(_05996_),
    .B(_06000_),
    .C(_06023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06025_));
 sky130_fd_sc_hd__or2_1 _12219_ (.A(_06024_),
    .B(_06025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06026_));
 sky130_fd_sc_hd__nand2_1 _12220_ (.A(_05983_),
    .B(_06005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06027_));
 sky130_fd_sc_hd__a21o_1 _12221_ (.A1(_05981_),
    .A2(_06004_),
    .B1(_06003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06028_));
 sky130_fd_sc_hd__o21a_1 _12222_ (.A1(_05967_),
    .A2(_06027_),
    .B1(_06028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06029_));
 sky130_fd_sc_hd__nor2_1 _12223_ (.A(_06026_),
    .B(_06029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06030_));
 sky130_fd_sc_hd__a211oi_1 _12224_ (.A1(_06026_),
    .A2(_06029_),
    .B1(_06030_),
    .C1(_05465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06031_));
 sky130_fd_sc_hd__a211o_1 _12225_ (.A1(\sha256cu.data_in_padd[26] ),
    .A2(_05667_),
    .B1(_06031_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06032_));
 sky130_fd_sc_hd__o211a_1 _12226_ (.A1(\sha256cu.iter_processing.w[26] ),
    .A2(_05894_),
    .B1(_06032_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00924_));
 sky130_fd_sc_hd__or2_1 _12227_ (.A(\sha256cu.msg_scheduler.mreg_9[27] ),
    .B(\sha256cu.msg_scheduler.mreg_0[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06033_));
 sky130_fd_sc_hd__nand2_1 _12228_ (.A(\sha256cu.msg_scheduler.mreg_9[27] ),
    .B(\sha256cu.msg_scheduler.mreg_0[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _12229_ (.A(_06033_),
    .B(_06034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06035_));
 sky130_fd_sc_hd__xnor2_1 _12230_ (.A(\sha256cu.msg_scheduler.mreg_1[13] ),
    .B(\sha256cu.msg_scheduler.mreg_1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06036_));
 sky130_fd_sc_hd__xnor2_1 _12231_ (.A(\sha256cu.msg_scheduler.mreg_1[30] ),
    .B(_06036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06037_));
 sky130_fd_sc_hd__xor2_1 _12232_ (.A(_06035_),
    .B(_06037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06038_));
 sky130_fd_sc_hd__a21boi_1 _12233_ (.A1(_06010_),
    .A2(_06014_),
    .B1_N(_06011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06039_));
 sky130_fd_sc_hd__nor2_1 _12234_ (.A(_06038_),
    .B(_06039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06040_));
 sky130_fd_sc_hd__and2_1 _12235_ (.A(_06038_),
    .B(_06039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06041_));
 sky130_fd_sc_hd__nor2_1 _12236_ (.A(_06040_),
    .B(_06041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06042_));
 sky130_fd_sc_hd__xor2_1 _12237_ (.A(\sha256cu.msg_scheduler.mreg_14[14] ),
    .B(\sha256cu.msg_scheduler.mreg_14[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06043_));
 sky130_fd_sc_hd__xnor2_1 _12238_ (.A(_06042_),
    .B(_06043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06044_));
 sky130_fd_sc_hd__nand3_1 _12239_ (.A(_06017_),
    .B(_06021_),
    .C(_06044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06045_));
 sky130_fd_sc_hd__inv_2 _12240_ (.A(_06045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06046_));
 sky130_fd_sc_hd__a21oi_1 _12241_ (.A1(_06017_),
    .A2(_06021_),
    .B1(_06044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06047_));
 sky130_fd_sc_hd__nor2_1 _12242_ (.A(_06046_),
    .B(_06047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06048_));
 sky130_fd_sc_hd__o21ai_1 _12243_ (.A1(_06024_),
    .A2(_06030_),
    .B1(_06048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06049_));
 sky130_fd_sc_hd__or3_1 _12244_ (.A(_06024_),
    .B(_06030_),
    .C(_06048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06050_));
 sky130_fd_sc_hd__a21o_1 _12245_ (.A1(\sha256cu.data_in_padd[27] ),
    .A2(_05447_),
    .B1(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06051_));
 sky130_fd_sc_hd__a31o_1 _12246_ (.A1(_05442_),
    .A2(_06049_),
    .A3(_06050_),
    .B1(_06051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06052_));
 sky130_fd_sc_hd__o211a_1 _12247_ (.A1(\sha256cu.iter_processing.w[27] ),
    .A2(_05894_),
    .B1(_06052_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00925_));
 sky130_fd_sc_hd__or3_1 _12248_ (.A(_06026_),
    .B(_06046_),
    .C(_06047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06053_));
 sky130_fd_sc_hd__a211o_1 _12249_ (.A1(_05963_),
    .A2(_05966_),
    .B1(_06027_),
    .C1(_06053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06054_));
 sky130_fd_sc_hd__a21oi_1 _12250_ (.A1(_06024_),
    .A2(_06045_),
    .B1(_06047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06055_));
 sky130_fd_sc_hd__o21a_1 _12251_ (.A1(_06028_),
    .A2(_06053_),
    .B1(_06055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06056_));
 sky130_fd_sc_hd__nand2_1 _12252_ (.A(\sha256cu.msg_scheduler.mreg_9[28] ),
    .B(\sha256cu.msg_scheduler.mreg_0[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06057_));
 sky130_fd_sc_hd__or2_1 _12253_ (.A(\sha256cu.msg_scheduler.mreg_9[28] ),
    .B(\sha256cu.msg_scheduler.mreg_0[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06058_));
 sky130_fd_sc_hd__nand2_1 _12254_ (.A(_06057_),
    .B(_06058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06059_));
 sky130_fd_sc_hd__xnor2_1 _12255_ (.A(\sha256cu.msg_scheduler.mreg_1[14] ),
    .B(\sha256cu.msg_scheduler.mreg_1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06060_));
 sky130_fd_sc_hd__xnor2_1 _12256_ (.A(\sha256cu.msg_scheduler.mreg_1[31] ),
    .B(_06060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06061_));
 sky130_fd_sc_hd__xor2_1 _12257_ (.A(_06059_),
    .B(_06061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06062_));
 sky130_fd_sc_hd__a21boi_1 _12258_ (.A1(_06033_),
    .A2(_06037_),
    .B1_N(_06034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06063_));
 sky130_fd_sc_hd__or2_2 _12259_ (.A(_06062_),
    .B(_06063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06064_));
 sky130_fd_sc_hd__nand2_1 _12260_ (.A(_06062_),
    .B(_06063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06065_));
 sky130_fd_sc_hd__and2_1 _12261_ (.A(_06064_),
    .B(_06065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06066_));
 sky130_fd_sc_hd__xor2_1 _12262_ (.A(\sha256cu.msg_scheduler.mreg_14[15] ),
    .B(\sha256cu.msg_scheduler.mreg_14[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06067_));
 sky130_fd_sc_hd__nand2_1 _12263_ (.A(_06066_),
    .B(_06067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06068_));
 sky130_fd_sc_hd__or2_1 _12264_ (.A(_06066_),
    .B(_06067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06069_));
 sky130_fd_sc_hd__nand2_1 _12265_ (.A(_06068_),
    .B(_06069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06070_));
 sky130_fd_sc_hd__a21oi_1 _12266_ (.A1(_06042_),
    .A2(_06043_),
    .B1(_06040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06071_));
 sky130_fd_sc_hd__nor2_2 _12267_ (.A(_06070_),
    .B(_06071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06072_));
 sky130_fd_sc_hd__and2_1 _12268_ (.A(_06070_),
    .B(_06071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06073_));
 sky130_fd_sc_hd__or2_1 _12269_ (.A(_06072_),
    .B(_06073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06074_));
 sky130_fd_sc_hd__a21oi_4 _12270_ (.A1(_06054_),
    .A2(_06056_),
    .B1(_06074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06075_));
 sky130_fd_sc_hd__and3_1 _12271_ (.A(_06074_),
    .B(_06054_),
    .C(_06056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06076_));
 sky130_fd_sc_hd__a21oi_1 _12272_ (.A1(\sha256cu.data_in_padd[28] ),
    .A2(_05433_),
    .B1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06077_));
 sky130_fd_sc_hd__o31ai_1 _12273_ (.A1(_05448_),
    .A2(_06075_),
    .A3(_06076_),
    .B1(_06077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06078_));
 sky130_fd_sc_hd__o211a_1 _12274_ (.A1(\sha256cu.iter_processing.w[28] ),
    .A2(_05894_),
    .B1(_06078_),
    .C1(_05866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00926_));
 sky130_fd_sc_hd__nand2_1 _12275_ (.A(\sha256cu.msg_scheduler.mreg_9[29] ),
    .B(\sha256cu.msg_scheduler.mreg_0[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06079_));
 sky130_fd_sc_hd__or2_1 _12276_ (.A(\sha256cu.msg_scheduler.mreg_9[29] ),
    .B(\sha256cu.msg_scheduler.mreg_0[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06080_));
 sky130_fd_sc_hd__nand2_1 _12277_ (.A(_06079_),
    .B(_06080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06081_));
 sky130_fd_sc_hd__xor2_1 _12278_ (.A(\sha256cu.msg_scheduler.mreg_1[15] ),
    .B(\sha256cu.msg_scheduler.mreg_1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06082_));
 sky130_fd_sc_hd__xor2_1 _12279_ (.A(_06081_),
    .B(_06082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06083_));
 sky130_fd_sc_hd__a21boi_1 _12280_ (.A1(_06058_),
    .A2(_06061_),
    .B1_N(_06057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06084_));
 sky130_fd_sc_hd__nor2_1 _12281_ (.A(_06083_),
    .B(_06084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06085_));
 sky130_fd_sc_hd__and2_1 _12282_ (.A(_06083_),
    .B(_06084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06086_));
 sky130_fd_sc_hd__nor2_2 _12283_ (.A(_06085_),
    .B(_06086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06087_));
 sky130_fd_sc_hd__xor2_2 _12284_ (.A(\sha256cu.msg_scheduler.mreg_14[16] ),
    .B(\sha256cu.msg_scheduler.mreg_14[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06088_));
 sky130_fd_sc_hd__xnor2_2 _12285_ (.A(_06087_),
    .B(_06088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06089_));
 sky130_fd_sc_hd__a21oi_2 _12286_ (.A1(_06064_),
    .A2(_06068_),
    .B1(_06089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06090_));
 sky130_fd_sc_hd__nand3_2 _12287_ (.A(_06064_),
    .B(_06068_),
    .C(_06089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06091_));
 sky130_fd_sc_hd__and2b_1 _12288_ (.A_N(_06090_),
    .B(_06091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06092_));
 sky130_fd_sc_hd__o21ai_1 _12289_ (.A1(_06072_),
    .A2(_06075_),
    .B1(_06092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06093_));
 sky130_fd_sc_hd__or3_1 _12290_ (.A(_06072_),
    .B(_06075_),
    .C(_06092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06094_));
 sky130_fd_sc_hd__a21o_1 _12291_ (.A1(\sha256cu.data_in_padd[29] ),
    .A2(_05447_),
    .B1(_04053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06095_));
 sky130_fd_sc_hd__a31o_1 _12292_ (.A1(_05442_),
    .A2(_06093_),
    .A3(_06094_),
    .B1(_06095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06096_));
 sky130_fd_sc_hd__o211a_1 _12293_ (.A1(\sha256cu.iter_processing.w[29] ),
    .A2(_05894_),
    .B1(_06096_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00927_));
 sky130_fd_sc_hd__or2_1 _12294_ (.A(\sha256cu.msg_scheduler.mreg_9[30] ),
    .B(\sha256cu.msg_scheduler.mreg_0[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06097_));
 sky130_fd_sc_hd__nand2_1 _12295_ (.A(\sha256cu.msg_scheduler.mreg_9[30] ),
    .B(\sha256cu.msg_scheduler.mreg_0[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_1 _12296_ (.A(_06097_),
    .B(_06098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06099_));
 sky130_fd_sc_hd__xor2_1 _12297_ (.A(\sha256cu.msg_scheduler.mreg_1[16] ),
    .B(\sha256cu.msg_scheduler.mreg_1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06100_));
 sky130_fd_sc_hd__xor2_1 _12298_ (.A(_06099_),
    .B(_06100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06101_));
 sky130_fd_sc_hd__a21boi_1 _12299_ (.A1(_06080_),
    .A2(_06082_),
    .B1_N(_06079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06102_));
 sky130_fd_sc_hd__xor2_1 _12300_ (.A(_06101_),
    .B(_06102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06103_));
 sky130_fd_sc_hd__xor2_1 _12301_ (.A(\sha256cu.msg_scheduler.mreg_14[17] ),
    .B(\sha256cu.msg_scheduler.mreg_14[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06104_));
 sky130_fd_sc_hd__nand2_1 _12302_ (.A(_06103_),
    .B(_06104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06105_));
 sky130_fd_sc_hd__or2_1 _12303_ (.A(_06103_),
    .B(_06104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06106_));
 sky130_fd_sc_hd__nand2_1 _12304_ (.A(_06105_),
    .B(_06106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06107_));
 sky130_fd_sc_hd__a21oi_1 _12305_ (.A1(_06087_),
    .A2(_06088_),
    .B1(_06085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06108_));
 sky130_fd_sc_hd__or2_1 _12306_ (.A(_06107_),
    .B(_06108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06109_));
 sky130_fd_sc_hd__nand2_1 _12307_ (.A(_06107_),
    .B(_06108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06110_));
 sky130_fd_sc_hd__and2_1 _12308_ (.A(_06109_),
    .B(_06110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06111_));
 sky130_fd_sc_hd__o311ai_4 _12309_ (.A1(_06072_),
    .A2(_06075_),
    .A3(_06090_),
    .B1(_06091_),
    .C1(_06111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06112_));
 sky130_fd_sc_hd__or2_1 _12310_ (.A(_06072_),
    .B(_06090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06113_));
 sky130_fd_sc_hd__a221o_1 _12311_ (.A1(_06075_),
    .A2(_06092_),
    .B1(_06113_),
    .B2(_06091_),
    .C1(_06111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06114_));
 sky130_fd_sc_hd__nand2_1 _12312_ (.A(_06112_),
    .B(_06114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06115_));
 sky130_fd_sc_hd__a21oi_1 _12313_ (.A1(\sha256cu.data_in_padd[30] ),
    .A2(_05433_),
    .B1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06116_));
 sky130_fd_sc_hd__o21ai_1 _12314_ (.A1(_05448_),
    .A2(_06115_),
    .B1(_06116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06117_));
 sky130_fd_sc_hd__o211a_1 _12315_ (.A1(\sha256cu.iter_processing.w[30] ),
    .A2(_05894_),
    .B1(_06117_),
    .C1(_01974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00928_));
 sky130_fd_sc_hd__o21a_1 _12316_ (.A1(_06101_),
    .A2(_06102_),
    .B1(_06105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06118_));
 sky130_fd_sc_hd__xnor2_1 _12317_ (.A(\sha256cu.msg_scheduler.mreg_14[18] ),
    .B(\sha256cu.msg_scheduler.mreg_14[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06119_));
 sky130_fd_sc_hd__xnor2_1 _12318_ (.A(\sha256cu.msg_scheduler.mreg_1[17] ),
    .B(_06119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06120_));
 sky130_fd_sc_hd__xor2_1 _12319_ (.A(\sha256cu.msg_scheduler.mreg_9[31] ),
    .B(\sha256cu.msg_scheduler.mreg_1[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06121_));
 sky130_fd_sc_hd__xnor2_1 _12320_ (.A(\sha256cu.msg_scheduler.mreg_0[31] ),
    .B(_06121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06122_));
 sky130_fd_sc_hd__xnor2_1 _12321_ (.A(_06120_),
    .B(_06122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06123_));
 sky130_fd_sc_hd__a21bo_1 _12322_ (.A1(_06097_),
    .A2(_06100_),
    .B1_N(_06098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06124_));
 sky130_fd_sc_hd__xnor2_1 _12323_ (.A(_06123_),
    .B(_06124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06125_));
 sky130_fd_sc_hd__xnor2_1 _12324_ (.A(_06118_),
    .B(_06125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06126_));
 sky130_fd_sc_hd__a21oi_1 _12325_ (.A1(_06109_),
    .A2(_06112_),
    .B1(_06126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06127_));
 sky130_fd_sc_hd__a31o_1 _12326_ (.A1(_06109_),
    .A2(_06112_),
    .A3(_06126_),
    .B1(_05465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06128_));
 sky130_fd_sc_hd__nor2_1 _12327_ (.A(_06127_),
    .B(_06128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06129_));
 sky130_fd_sc_hd__a21o_1 _12328_ (.A1(\sha256cu.data_in_padd[31] ),
    .A2(_05448_),
    .B1(_05463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06130_));
 sky130_fd_sc_hd__o221a_1 _12329_ (.A1(\sha256cu.iter_processing.w[31] ),
    .A2(_04044_),
    .B1(_06129_),
    .B2(_06130_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00929_));
 sky130_fd_sc_hd__and2_1 _12330_ (.A(_03288_),
    .B(_01949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06131_));
 sky130_fd_sc_hd__clkbuf_1 _12331_ (.A(_06131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00930_));
 sky130_fd_sc_hd__and3_1 _12332_ (.A(\sha256cu.m_pad_pars.add_512_block[1] ),
    .B(_01939_),
    .C(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06132_));
 sky130_fd_sc_hd__a21o_1 _12333_ (.A1(_01939_),
    .A2(_01947_),
    .B1(\sha256cu.m_pad_pars.add_512_block[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06133_));
 sky130_fd_sc_hd__and3b_1 _12334_ (.A_N(_06132_),
    .B(_01983_),
    .C(_06133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06134_));
 sky130_fd_sc_hd__clkbuf_1 _12335_ (.A(_06134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00931_));
 sky130_fd_sc_hd__o21ai_1 _12336_ (.A1(\sha256cu.m_pad_pars.add_512_block[2] ),
    .A2(_06132_),
    .B1(_03288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06135_));
 sky130_fd_sc_hd__a21oi_1 _12337_ (.A1(\sha256cu.m_pad_pars.add_512_block[2] ),
    .A2(_06132_),
    .B1(_06135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00932_));
 sky130_fd_sc_hd__and2_1 _12338_ (.A(_01947_),
    .B(_04777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06136_));
 sky130_fd_sc_hd__a21o_1 _12339_ (.A1(\sha256cu.m_pad_pars.add_512_block[2] ),
    .A2(_06132_),
    .B1(\sha256cu.m_pad_pars.add_512_block[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06137_));
 sky130_fd_sc_hd__and3b_1 _12340_ (.A_N(_06136_),
    .B(_01983_),
    .C(_06137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06138_));
 sky130_fd_sc_hd__clkbuf_1 _12341_ (.A(_06138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00933_));
 sky130_fd_sc_hd__or2_1 _12342_ (.A(\sha256cu.m_pad_pars.add_512_block[4] ),
    .B(_06136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06139_));
 sky130_fd_sc_hd__nand2_1 _12343_ (.A(\sha256cu.m_pad_pars.add_512_block[4] ),
    .B(_06136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06140_));
 sky130_fd_sc_hd__and3_1 _12344_ (.A(_01973_),
    .B(_06139_),
    .C(_06140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06141_));
 sky130_fd_sc_hd__clkbuf_1 _12345_ (.A(_06141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00934_));
 sky130_fd_sc_hd__and3_1 _12346_ (.A(\sha256cu.byte_rdy ),
    .B(_01914_),
    .C(_04777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06142_));
 sky130_fd_sc_hd__a211oi_1 _12347_ (.A1(_04743_),
    .A2(_06140_),
    .B1(_06142_),
    .C1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00935_));
 sky130_fd_sc_hd__a21o_1 _12348_ (.A1(\sha256cu.m_pad_pars.add_512_block[6] ),
    .A2(_06142_),
    .B1(_02002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06143_));
 sky130_fd_sc_hd__o21ba_1 _12349_ (.A1(\sha256cu.m_pad_pars.add_512_block[6] ),
    .A2(_06142_),
    .B1_N(_06143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00936_));
 sky130_fd_sc_hd__or3_2 _12350_ (.A(_01986_),
    .B(_05264_),
    .C(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06144_));
 sky130_fd_sc_hd__and2_1 _12351_ (.A(\sha256cu.m_pad_pars.block_512[0][0] ),
    .B(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06145_));
 sky130_fd_sc_hd__clkbuf_1 _12352_ (.A(_06145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00937_));
 sky130_fd_sc_hd__and2_1 _12353_ (.A(\sha256cu.m_pad_pars.block_512[0][1] ),
    .B(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06146_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_06146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00938_));
 sky130_fd_sc_hd__and2_1 _12355_ (.A(\sha256cu.m_pad_pars.block_512[0][2] ),
    .B(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06147_));
 sky130_fd_sc_hd__clkbuf_1 _12356_ (.A(_06147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00939_));
 sky130_fd_sc_hd__and2_1 _12357_ (.A(\sha256cu.m_pad_pars.block_512[0][3] ),
    .B(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_1 _12358_ (.A(_06148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00940_));
 sky130_fd_sc_hd__and2_1 _12359_ (.A(\sha256cu.m_pad_pars.block_512[0][4] ),
    .B(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06149_));
 sky130_fd_sc_hd__clkbuf_1 _12360_ (.A(_06149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00941_));
 sky130_fd_sc_hd__and2_1 _12361_ (.A(\sha256cu.m_pad_pars.block_512[0][5] ),
    .B(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_1 _12362_ (.A(_06150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00942_));
 sky130_fd_sc_hd__and2_1 _12363_ (.A(\sha256cu.m_pad_pars.block_512[0][6] ),
    .B(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _12364_ (.A(_06151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00943_));
 sky130_fd_sc_hd__a31o_1 _12365_ (.A1(_01984_),
    .A2(_01942_),
    .A3(_04775_),
    .B1(\sha256cu.m_pad_pars.block_512[0][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00944_));
 sky130_fd_sc_hd__nand2_2 _12366_ (.A(_01965_),
    .B(_05244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06152_));
 sky130_fd_sc_hd__and2_1 _12367_ (.A(\sha256cu.m_pad_pars.block_512[1][0] ),
    .B(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06153_));
 sky130_fd_sc_hd__clkbuf_1 _12368_ (.A(_06153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00945_));
 sky130_fd_sc_hd__and2_1 _12369_ (.A(\sha256cu.m_pad_pars.block_512[1][1] ),
    .B(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_1 _12370_ (.A(_06154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00946_));
 sky130_fd_sc_hd__and2_1 _12371_ (.A(\sha256cu.m_pad_pars.block_512[1][2] ),
    .B(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06155_));
 sky130_fd_sc_hd__clkbuf_1 _12372_ (.A(_06155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00947_));
 sky130_fd_sc_hd__and2_1 _12373_ (.A(\sha256cu.m_pad_pars.block_512[1][3] ),
    .B(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06156_));
 sky130_fd_sc_hd__clkbuf_1 _12374_ (.A(_06156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00948_));
 sky130_fd_sc_hd__and2_1 _12375_ (.A(\sha256cu.m_pad_pars.block_512[1][4] ),
    .B(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_1 _12376_ (.A(_06157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00949_));
 sky130_fd_sc_hd__and2_1 _12377_ (.A(\sha256cu.m_pad_pars.block_512[1][5] ),
    .B(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06158_));
 sky130_fd_sc_hd__clkbuf_1 _12378_ (.A(_06158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00950_));
 sky130_fd_sc_hd__and2_1 _12379_ (.A(\sha256cu.m_pad_pars.block_512[1][6] ),
    .B(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_1 _12380_ (.A(_06159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00951_));
 sky130_fd_sc_hd__a21o_1 _12381_ (.A1(_02000_),
    .A2(_05244_),
    .B1(\sha256cu.m_pad_pars.block_512[1][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00952_));
 sky130_fd_sc_hd__nand2_2 _12382_ (.A(_01965_),
    .B(_04998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06160_));
 sky130_fd_sc_hd__and2_1 _12383_ (.A(\sha256cu.m_pad_pars.block_512[2][0] ),
    .B(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_1 _12384_ (.A(_06161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00953_));
 sky130_fd_sc_hd__and2_1 _12385_ (.A(\sha256cu.m_pad_pars.block_512[2][1] ),
    .B(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_1 _12386_ (.A(_06162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00954_));
 sky130_fd_sc_hd__and2_1 _12387_ (.A(\sha256cu.m_pad_pars.block_512[2][2] ),
    .B(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06163_));
 sky130_fd_sc_hd__clkbuf_1 _12388_ (.A(_06163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00955_));
 sky130_fd_sc_hd__and2_1 _12389_ (.A(\sha256cu.m_pad_pars.block_512[2][3] ),
    .B(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06164_));
 sky130_fd_sc_hd__clkbuf_1 _12390_ (.A(_06164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00956_));
 sky130_fd_sc_hd__and2_1 _12391_ (.A(\sha256cu.m_pad_pars.block_512[2][4] ),
    .B(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06165_));
 sky130_fd_sc_hd__clkbuf_1 _12392_ (.A(_06165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00957_));
 sky130_fd_sc_hd__and2_1 _12393_ (.A(\sha256cu.m_pad_pars.block_512[2][5] ),
    .B(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06166_));
 sky130_fd_sc_hd__clkbuf_1 _12394_ (.A(_06166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00958_));
 sky130_fd_sc_hd__and2_1 _12395_ (.A(\sha256cu.m_pad_pars.block_512[2][6] ),
    .B(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06167_));
 sky130_fd_sc_hd__clkbuf_1 _12396_ (.A(_06167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00959_));
 sky130_fd_sc_hd__nor2_1 _12397_ (.A(_03288_),
    .B(\sha256cu.m_pad_pars.block_512[2][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06168_));
 sky130_fd_sc_hd__a21oi_1 _12398_ (.A1(_01966_),
    .A2(_05119_),
    .B1(_06168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00960_));
 sky130_fd_sc_hd__nand2_2 _12399_ (.A(_01965_),
    .B(_04763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06169_));
 sky130_fd_sc_hd__and2_1 _12400_ (.A(\sha256cu.m_pad_pars.block_512[3][0] ),
    .B(_06169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _12401_ (.A(_06170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00961_));
 sky130_fd_sc_hd__and2_1 _12402_ (.A(\sha256cu.m_pad_pars.block_512[3][1] ),
    .B(_06169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06171_));
 sky130_fd_sc_hd__clkbuf_1 _12403_ (.A(_06171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00962_));
 sky130_fd_sc_hd__and2_1 _12404_ (.A(\sha256cu.m_pad_pars.block_512[3][2] ),
    .B(_06169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _12405_ (.A(_06172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00963_));
 sky130_fd_sc_hd__and2_1 _12406_ (.A(\sha256cu.m_pad_pars.block_512[3][3] ),
    .B(_06169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06173_));
 sky130_fd_sc_hd__clkbuf_1 _12407_ (.A(_06173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00964_));
 sky130_fd_sc_hd__and2_1 _12408_ (.A(\sha256cu.m_pad_pars.block_512[3][4] ),
    .B(_06169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_1 _12409_ (.A(_06174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00965_));
 sky130_fd_sc_hd__and2_1 _12410_ (.A(\sha256cu.m_pad_pars.block_512[3][5] ),
    .B(_06169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_1 _12411_ (.A(_06175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00966_));
 sky130_fd_sc_hd__and2_1 _12412_ (.A(\sha256cu.m_pad_pars.block_512[3][6] ),
    .B(_06169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06176_));
 sky130_fd_sc_hd__clkbuf_1 _12413_ (.A(_06176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(\sha256cu.m_pad_pars.block_512[3][7] ),
    .A1(_04935_),
    .S(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06177_));
 sky130_fd_sc_hd__clkbuf_1 _12415_ (.A(_06177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00968_));
 sky130_fd_sc_hd__or2_2 _12416_ (.A(_01912_),
    .B(_05312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06178_));
 sky130_fd_sc_hd__and2_1 _12417_ (.A(\sha256cu.m_pad_pars.block_512[4][0] ),
    .B(_06178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06179_));
 sky130_fd_sc_hd__clkbuf_1 _12418_ (.A(_06179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00969_));
 sky130_fd_sc_hd__and2_1 _12419_ (.A(\sha256cu.m_pad_pars.block_512[4][1] ),
    .B(_06178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06180_));
 sky130_fd_sc_hd__clkbuf_1 _12420_ (.A(_06180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00970_));
 sky130_fd_sc_hd__and2_1 _12421_ (.A(\sha256cu.m_pad_pars.block_512[4][2] ),
    .B(_06178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06181_));
 sky130_fd_sc_hd__clkbuf_1 _12422_ (.A(_06181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00971_));
 sky130_fd_sc_hd__and2_1 _12423_ (.A(\sha256cu.m_pad_pars.block_512[4][3] ),
    .B(_06178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06182_));
 sky130_fd_sc_hd__clkbuf_1 _12424_ (.A(_06182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00972_));
 sky130_fd_sc_hd__and2_1 _12425_ (.A(\sha256cu.m_pad_pars.block_512[4][4] ),
    .B(_06178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06183_));
 sky130_fd_sc_hd__clkbuf_1 _12426_ (.A(_06183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00973_));
 sky130_fd_sc_hd__and2_1 _12427_ (.A(\sha256cu.m_pad_pars.block_512[4][5] ),
    .B(_06178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06184_));
 sky130_fd_sc_hd__clkbuf_1 _12428_ (.A(_06184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00974_));
 sky130_fd_sc_hd__and2_1 _12429_ (.A(\sha256cu.m_pad_pars.block_512[4][6] ),
    .B(_06178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06185_));
 sky130_fd_sc_hd__clkbuf_1 _12430_ (.A(_06185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _12431_ (.A0(\sha256cu.m_pad_pars.block_512[4][7] ),
    .A1(_05411_),
    .S(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06186_));
 sky130_fd_sc_hd__clkbuf_1 _12432_ (.A(_06186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00976_));
 sky130_fd_sc_hd__or3_2 _12433_ (.A(_01986_),
    .B(_04933_),
    .C(_05159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06187_));
 sky130_fd_sc_hd__and2_1 _12434_ (.A(\sha256cu.m_pad_pars.block_512[5][0] ),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06188_));
 sky130_fd_sc_hd__clkbuf_1 _12435_ (.A(_06188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00977_));
 sky130_fd_sc_hd__and2_1 _12436_ (.A(\sha256cu.m_pad_pars.block_512[5][1] ),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06189_));
 sky130_fd_sc_hd__clkbuf_1 _12437_ (.A(_06189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00978_));
 sky130_fd_sc_hd__and2_1 _12438_ (.A(\sha256cu.m_pad_pars.block_512[5][2] ),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06190_));
 sky130_fd_sc_hd__clkbuf_1 _12439_ (.A(_06190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00979_));
 sky130_fd_sc_hd__and2_1 _12440_ (.A(\sha256cu.m_pad_pars.block_512[5][3] ),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06191_));
 sky130_fd_sc_hd__clkbuf_1 _12441_ (.A(_06191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00980_));
 sky130_fd_sc_hd__and2_1 _12442_ (.A(\sha256cu.m_pad_pars.block_512[5][4] ),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_1 _12443_ (.A(_06192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00981_));
 sky130_fd_sc_hd__and2_1 _12444_ (.A(\sha256cu.m_pad_pars.block_512[5][5] ),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06193_));
 sky130_fd_sc_hd__clkbuf_1 _12445_ (.A(_06193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00982_));
 sky130_fd_sc_hd__and2_1 _12446_ (.A(\sha256cu.m_pad_pars.block_512[5][6] ),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06194_));
 sky130_fd_sc_hd__clkbuf_1 _12447_ (.A(_06194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _12448_ (.A0(\sha256cu.m_pad_pars.block_512[5][7] ),
    .A1(_05238_),
    .S(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06195_));
 sky130_fd_sc_hd__clkbuf_1 _12449_ (.A(_06195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00984_));
 sky130_fd_sc_hd__nand2_2 _12450_ (.A(_01965_),
    .B(_04956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06196_));
 sky130_fd_sc_hd__and2_1 _12451_ (.A(\sha256cu.m_pad_pars.block_512[6][0] ),
    .B(_06196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06197_));
 sky130_fd_sc_hd__clkbuf_1 _12452_ (.A(_06197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00985_));
 sky130_fd_sc_hd__and2_1 _12453_ (.A(\sha256cu.m_pad_pars.block_512[6][1] ),
    .B(_06196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_06198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00986_));
 sky130_fd_sc_hd__and2_1 _12455_ (.A(\sha256cu.m_pad_pars.block_512[6][2] ),
    .B(_06196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06199_));
 sky130_fd_sc_hd__clkbuf_1 _12456_ (.A(_06199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00987_));
 sky130_fd_sc_hd__and2_1 _12457_ (.A(\sha256cu.m_pad_pars.block_512[6][3] ),
    .B(_06196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_1 _12458_ (.A(_06200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00988_));
 sky130_fd_sc_hd__and2_1 _12459_ (.A(\sha256cu.m_pad_pars.block_512[6][4] ),
    .B(_06196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06201_));
 sky130_fd_sc_hd__clkbuf_1 _12460_ (.A(_06201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00989_));
 sky130_fd_sc_hd__and2_1 _12461_ (.A(\sha256cu.m_pad_pars.block_512[6][5] ),
    .B(_06196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_1 _12462_ (.A(_06202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00990_));
 sky130_fd_sc_hd__and2_1 _12463_ (.A(\sha256cu.m_pad_pars.block_512[6][6] ),
    .B(_06196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06203_));
 sky130_fd_sc_hd__clkbuf_1 _12464_ (.A(_06203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(\sha256cu.m_pad_pars.block_512[6][7] ),
    .A1(_05099_),
    .S(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_1 _12466_ (.A(_06204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00992_));
 sky130_fd_sc_hd__or2_2 _12467_ (.A(_01912_),
    .B(_04773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06205_));
 sky130_fd_sc_hd__and2_1 _12468_ (.A(\sha256cu.m_pad_pars.block_512[7][0] ),
    .B(_06205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_1 _12469_ (.A(_06206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00993_));
 sky130_fd_sc_hd__and2_1 _12470_ (.A(\sha256cu.m_pad_pars.block_512[7][1] ),
    .B(_06205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_1 _12471_ (.A(_06207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00994_));
 sky130_fd_sc_hd__and2_1 _12472_ (.A(\sha256cu.m_pad_pars.block_512[7][2] ),
    .B(_06205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06208_));
 sky130_fd_sc_hd__clkbuf_1 _12473_ (.A(_06208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00995_));
 sky130_fd_sc_hd__and2_1 _12474_ (.A(\sha256cu.m_pad_pars.block_512[7][3] ),
    .B(_06205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06209_));
 sky130_fd_sc_hd__clkbuf_1 _12475_ (.A(_06209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00996_));
 sky130_fd_sc_hd__and2_1 _12476_ (.A(\sha256cu.m_pad_pars.block_512[7][4] ),
    .B(_06205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_1 _12477_ (.A(_06210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00997_));
 sky130_fd_sc_hd__and2_1 _12478_ (.A(\sha256cu.m_pad_pars.block_512[7][5] ),
    .B(_06205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06211_));
 sky130_fd_sc_hd__clkbuf_1 _12479_ (.A(_06211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00998_));
 sky130_fd_sc_hd__and2_1 _12480_ (.A(\sha256cu.m_pad_pars.block_512[7][6] ),
    .B(_06205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06212_));
 sky130_fd_sc_hd__clkbuf_1 _12481_ (.A(_06212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _12482_ (.A0(\sha256cu.m_pad_pars.block_512[7][7] ),
    .A1(_04923_),
    .S(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06213_));
 sky130_fd_sc_hd__clkbuf_1 _12483_ (.A(_06213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01000_));
 sky130_fd_sc_hd__nand2_2 _12484_ (.A(_01965_),
    .B(_05317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06214_));
 sky130_fd_sc_hd__and2_1 _12485_ (.A(\sha256cu.m_pad_pars.block_512[8][0] ),
    .B(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06215_));
 sky130_fd_sc_hd__clkbuf_1 _12486_ (.A(_06215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01001_));
 sky130_fd_sc_hd__and2_1 _12487_ (.A(\sha256cu.m_pad_pars.block_512[8][1] ),
    .B(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06216_));
 sky130_fd_sc_hd__clkbuf_1 _12488_ (.A(_06216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01002_));
 sky130_fd_sc_hd__and2_1 _12489_ (.A(\sha256cu.m_pad_pars.block_512[8][2] ),
    .B(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06217_));
 sky130_fd_sc_hd__clkbuf_1 _12490_ (.A(_06217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01003_));
 sky130_fd_sc_hd__and2_1 _12491_ (.A(\sha256cu.m_pad_pars.block_512[8][3] ),
    .B(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06218_));
 sky130_fd_sc_hd__clkbuf_1 _12492_ (.A(_06218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01004_));
 sky130_fd_sc_hd__and2_1 _12493_ (.A(\sha256cu.m_pad_pars.block_512[8][4] ),
    .B(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06219_));
 sky130_fd_sc_hd__clkbuf_1 _12494_ (.A(_06219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01005_));
 sky130_fd_sc_hd__and2_1 _12495_ (.A(\sha256cu.m_pad_pars.block_512[8][5] ),
    .B(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06220_));
 sky130_fd_sc_hd__clkbuf_1 _12496_ (.A(_06220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01006_));
 sky130_fd_sc_hd__and2_1 _12497_ (.A(\sha256cu.m_pad_pars.block_512[8][6] ),
    .B(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06221_));
 sky130_fd_sc_hd__clkbuf_1 _12498_ (.A(_06221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(\sha256cu.m_pad_pars.block_512[8][7] ),
    .A1(_05424_),
    .S(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_1 _12500_ (.A(_06222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01008_));
 sky130_fd_sc_hd__or3_2 _12501_ (.A(_01986_),
    .B(_04933_),
    .C(_05130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06223_));
 sky130_fd_sc_hd__and2_1 _12502_ (.A(\sha256cu.m_pad_pars.block_512[9][0] ),
    .B(_06223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06224_));
 sky130_fd_sc_hd__clkbuf_1 _12503_ (.A(_06224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01009_));
 sky130_fd_sc_hd__and2_1 _12504_ (.A(\sha256cu.m_pad_pars.block_512[9][1] ),
    .B(_06223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06225_));
 sky130_fd_sc_hd__clkbuf_1 _12505_ (.A(_06225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01010_));
 sky130_fd_sc_hd__and2_1 _12506_ (.A(\sha256cu.m_pad_pars.block_512[9][2] ),
    .B(_06223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_1 _12507_ (.A(_06226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01011_));
 sky130_fd_sc_hd__and2_1 _12508_ (.A(\sha256cu.m_pad_pars.block_512[9][3] ),
    .B(_06223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06227_));
 sky130_fd_sc_hd__clkbuf_1 _12509_ (.A(_06227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01012_));
 sky130_fd_sc_hd__and2_1 _12510_ (.A(\sha256cu.m_pad_pars.block_512[9][4] ),
    .B(_06223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06228_));
 sky130_fd_sc_hd__clkbuf_1 _12511_ (.A(_06228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01013_));
 sky130_fd_sc_hd__and2_1 _12512_ (.A(\sha256cu.m_pad_pars.block_512[9][5] ),
    .B(_06223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06229_));
 sky130_fd_sc_hd__clkbuf_1 _12513_ (.A(_06229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01014_));
 sky130_fd_sc_hd__and2_1 _12514_ (.A(\sha256cu.m_pad_pars.block_512[9][6] ),
    .B(_06223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06230_));
 sky130_fd_sc_hd__clkbuf_1 _12515_ (.A(_06230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(\sha256cu.m_pad_pars.block_512[9][7] ),
    .A1(_05260_),
    .S(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06231_));
 sky130_fd_sc_hd__clkbuf_1 _12517_ (.A(_06231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01016_));
 sky130_fd_sc_hd__nand2_2 _12518_ (.A(_01965_),
    .B(_04962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06232_));
 sky130_fd_sc_hd__and2_1 _12519_ (.A(\sha256cu.m_pad_pars.block_512[10][0] ),
    .B(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_1 _12520_ (.A(_06233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01017_));
 sky130_fd_sc_hd__and2_1 _12521_ (.A(\sha256cu.m_pad_pars.block_512[10][1] ),
    .B(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06234_));
 sky130_fd_sc_hd__clkbuf_1 _12522_ (.A(_06234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01018_));
 sky130_fd_sc_hd__and2_1 _12523_ (.A(\sha256cu.m_pad_pars.block_512[10][2] ),
    .B(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06235_));
 sky130_fd_sc_hd__clkbuf_1 _12524_ (.A(_06235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01019_));
 sky130_fd_sc_hd__and2_1 _12525_ (.A(\sha256cu.m_pad_pars.block_512[10][3] ),
    .B(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06236_));
 sky130_fd_sc_hd__clkbuf_1 _12526_ (.A(_06236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01020_));
 sky130_fd_sc_hd__and2_1 _12527_ (.A(\sha256cu.m_pad_pars.block_512[10][4] ),
    .B(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06237_));
 sky130_fd_sc_hd__clkbuf_1 _12528_ (.A(_06237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01021_));
 sky130_fd_sc_hd__and2_1 _12529_ (.A(\sha256cu.m_pad_pars.block_512[10][5] ),
    .B(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_1 _12530_ (.A(_06238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01022_));
 sky130_fd_sc_hd__and2_1 _12531_ (.A(\sha256cu.m_pad_pars.block_512[10][6] ),
    .B(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_1 _12532_ (.A(_06239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01023_));
 sky130_fd_sc_hd__o211a_1 _12533_ (.A1(\sha256cu.m_pad_pars.block_512[10][7] ),
    .A2(_05090_),
    .B1(_05091_),
    .C1(_01975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06240_));
 sky130_fd_sc_hd__a21o_1 _12534_ (.A1(_02068_),
    .A2(\sha256cu.m_pad_pars.block_512[10][7] ),
    .B1(_06240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01024_));
 sky130_fd_sc_hd__nand2_2 _12535_ (.A(_01965_),
    .B(_04789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06241_));
 sky130_fd_sc_hd__and2_1 _12536_ (.A(\sha256cu.m_pad_pars.block_512[11][0] ),
    .B(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06242_));
 sky130_fd_sc_hd__clkbuf_1 _12537_ (.A(_06242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01025_));
 sky130_fd_sc_hd__and2_1 _12538_ (.A(\sha256cu.m_pad_pars.block_512[11][1] ),
    .B(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _12539_ (.A(_06243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01026_));
 sky130_fd_sc_hd__and2_1 _12540_ (.A(\sha256cu.m_pad_pars.block_512[11][2] ),
    .B(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_1 _12541_ (.A(_06244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01027_));
 sky130_fd_sc_hd__and2_1 _12542_ (.A(\sha256cu.m_pad_pars.block_512[11][3] ),
    .B(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_1 _12543_ (.A(_06245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01028_));
 sky130_fd_sc_hd__and2_1 _12544_ (.A(\sha256cu.m_pad_pars.block_512[11][4] ),
    .B(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_1 _12545_ (.A(_06246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01029_));
 sky130_fd_sc_hd__and2_1 _12546_ (.A(\sha256cu.m_pad_pars.block_512[11][5] ),
    .B(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06247_));
 sky130_fd_sc_hd__clkbuf_1 _12547_ (.A(_06247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01030_));
 sky130_fd_sc_hd__and2_1 _12548_ (.A(\sha256cu.m_pad_pars.block_512[11][6] ),
    .B(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _12549_ (.A(_06248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01031_));
 sky130_fd_sc_hd__buf_4 _12550_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06249_));
 sky130_fd_sc_hd__mux2_1 _12551_ (.A0(\sha256cu.m_pad_pars.block_512[11][7] ),
    .A1(_04946_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_1 _12552_ (.A(_06250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01032_));
 sky130_fd_sc_hd__buf_4 _12553_ (.A(_01911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06251_));
 sky130_fd_sc_hd__or3_2 _12554_ (.A(_06251_),
    .B(_04933_),
    .C(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06252_));
 sky130_fd_sc_hd__and2_1 _12555_ (.A(\sha256cu.m_pad_pars.block_512[12][0] ),
    .B(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06253_));
 sky130_fd_sc_hd__clkbuf_1 _12556_ (.A(_06253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01033_));
 sky130_fd_sc_hd__and2_1 _12557_ (.A(\sha256cu.m_pad_pars.block_512[12][1] ),
    .B(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06254_));
 sky130_fd_sc_hd__clkbuf_1 _12558_ (.A(_06254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01034_));
 sky130_fd_sc_hd__and2_1 _12559_ (.A(\sha256cu.m_pad_pars.block_512[12][2] ),
    .B(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06255_));
 sky130_fd_sc_hd__clkbuf_1 _12560_ (.A(_06255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01035_));
 sky130_fd_sc_hd__and2_1 _12561_ (.A(\sha256cu.m_pad_pars.block_512[12][3] ),
    .B(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06256_));
 sky130_fd_sc_hd__clkbuf_1 _12562_ (.A(_06256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01036_));
 sky130_fd_sc_hd__and2_1 _12563_ (.A(\sha256cu.m_pad_pars.block_512[12][4] ),
    .B(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06257_));
 sky130_fd_sc_hd__clkbuf_1 _12564_ (.A(_06257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01037_));
 sky130_fd_sc_hd__and2_1 _12565_ (.A(\sha256cu.m_pad_pars.block_512[12][5] ),
    .B(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06258_));
 sky130_fd_sc_hd__clkbuf_1 _12566_ (.A(_06258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01038_));
 sky130_fd_sc_hd__and2_1 _12567_ (.A(\sha256cu.m_pad_pars.block_512[12][6] ),
    .B(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06259_));
 sky130_fd_sc_hd__clkbuf_1 _12568_ (.A(_06259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _12569_ (.A0(\sha256cu.m_pad_pars.block_512[12][7] ),
    .A1(_05407_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_1 _12570_ (.A(_06260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01040_));
 sky130_fd_sc_hd__or3_2 _12571_ (.A(_06251_),
    .B(_04933_),
    .C(_05124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06261_));
 sky130_fd_sc_hd__and2_1 _12572_ (.A(\sha256cu.m_pad_pars.block_512[13][0] ),
    .B(_06261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06262_));
 sky130_fd_sc_hd__clkbuf_1 _12573_ (.A(_06262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01041_));
 sky130_fd_sc_hd__and2_1 _12574_ (.A(\sha256cu.m_pad_pars.block_512[13][1] ),
    .B(_06261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_1 _12575_ (.A(_06263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01042_));
 sky130_fd_sc_hd__and2_1 _12576_ (.A(\sha256cu.m_pad_pars.block_512[13][2] ),
    .B(_06261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06264_));
 sky130_fd_sc_hd__clkbuf_1 _12577_ (.A(_06264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01043_));
 sky130_fd_sc_hd__and2_1 _12578_ (.A(\sha256cu.m_pad_pars.block_512[13][3] ),
    .B(_06261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06265_));
 sky130_fd_sc_hd__clkbuf_1 _12579_ (.A(_06265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01044_));
 sky130_fd_sc_hd__and2_1 _12580_ (.A(\sha256cu.m_pad_pars.block_512[13][4] ),
    .B(_06261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06266_));
 sky130_fd_sc_hd__clkbuf_1 _12581_ (.A(_06266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01045_));
 sky130_fd_sc_hd__and2_1 _12582_ (.A(\sha256cu.m_pad_pars.block_512[13][5] ),
    .B(_06261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06267_));
 sky130_fd_sc_hd__clkbuf_1 _12583_ (.A(_06267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01046_));
 sky130_fd_sc_hd__and2_1 _12584_ (.A(\sha256cu.m_pad_pars.block_512[13][6] ),
    .B(_06261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06268_));
 sky130_fd_sc_hd__clkbuf_1 _12585_ (.A(_06268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _12586_ (.A0(\sha256cu.m_pad_pars.block_512[13][7] ),
    .A1(_05258_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06269_));
 sky130_fd_sc_hd__clkbuf_1 _12587_ (.A(_06269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01048_));
 sky130_fd_sc_hd__buf_6 _12588_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06270_));
 sky130_fd_sc_hd__nand2_2 _12589_ (.A(_06270_),
    .B(_04988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06271_));
 sky130_fd_sc_hd__and2_1 _12590_ (.A(\sha256cu.m_pad_pars.block_512[14][0] ),
    .B(_06271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06272_));
 sky130_fd_sc_hd__clkbuf_1 _12591_ (.A(_06272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01049_));
 sky130_fd_sc_hd__and2_1 _12592_ (.A(\sha256cu.m_pad_pars.block_512[14][1] ),
    .B(_06271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06273_));
 sky130_fd_sc_hd__clkbuf_1 _12593_ (.A(_06273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01050_));
 sky130_fd_sc_hd__and2_1 _12594_ (.A(\sha256cu.m_pad_pars.block_512[14][2] ),
    .B(_06271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06274_));
 sky130_fd_sc_hd__clkbuf_1 _12595_ (.A(_06274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01051_));
 sky130_fd_sc_hd__and2_1 _12596_ (.A(\sha256cu.m_pad_pars.block_512[14][3] ),
    .B(_06271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_1 _12597_ (.A(_06275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01052_));
 sky130_fd_sc_hd__and2_1 _12598_ (.A(\sha256cu.m_pad_pars.block_512[14][4] ),
    .B(_06271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06276_));
 sky130_fd_sc_hd__clkbuf_1 _12599_ (.A(_06276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01053_));
 sky130_fd_sc_hd__and2_1 _12600_ (.A(\sha256cu.m_pad_pars.block_512[14][5] ),
    .B(_06271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06277_));
 sky130_fd_sc_hd__clkbuf_1 _12601_ (.A(_06277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01054_));
 sky130_fd_sc_hd__and2_1 _12602_ (.A(\sha256cu.m_pad_pars.block_512[14][6] ),
    .B(_06271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06278_));
 sky130_fd_sc_hd__clkbuf_1 _12603_ (.A(_06278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(\sha256cu.m_pad_pars.block_512[14][7] ),
    .A1(_05097_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06279_));
 sky130_fd_sc_hd__clkbuf_1 _12605_ (.A(_06279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01056_));
 sky130_fd_sc_hd__a21o_2 _12606_ (.A1(_04778_),
    .A2(_04780_),
    .B1(_01912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06280_));
 sky130_fd_sc_hd__and2_1 _12607_ (.A(\sha256cu.m_pad_pars.block_512[15][0] ),
    .B(_06280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_1 _12608_ (.A(_06281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01057_));
 sky130_fd_sc_hd__and2_1 _12609_ (.A(\sha256cu.m_pad_pars.block_512[15][1] ),
    .B(_06280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_1 _12610_ (.A(_06282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01058_));
 sky130_fd_sc_hd__and2_1 _12611_ (.A(\sha256cu.m_pad_pars.block_512[15][2] ),
    .B(_06280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06283_));
 sky130_fd_sc_hd__clkbuf_1 _12612_ (.A(_06283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01059_));
 sky130_fd_sc_hd__and2_1 _12613_ (.A(\sha256cu.m_pad_pars.block_512[15][3] ),
    .B(_06280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06284_));
 sky130_fd_sc_hd__clkbuf_1 _12614_ (.A(_06284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01060_));
 sky130_fd_sc_hd__and2_1 _12615_ (.A(\sha256cu.m_pad_pars.block_512[15][4] ),
    .B(_06280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06285_));
 sky130_fd_sc_hd__clkbuf_1 _12616_ (.A(_06285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01061_));
 sky130_fd_sc_hd__and2_1 _12617_ (.A(\sha256cu.m_pad_pars.block_512[15][5] ),
    .B(_06280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06286_));
 sky130_fd_sc_hd__clkbuf_1 _12618_ (.A(_06286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01062_));
 sky130_fd_sc_hd__and2_1 _12619_ (.A(\sha256cu.m_pad_pars.block_512[15][6] ),
    .B(_06280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06287_));
 sky130_fd_sc_hd__clkbuf_1 _12620_ (.A(_06287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01063_));
 sky130_fd_sc_hd__nor2_1 _12621_ (.A(_03288_),
    .B(\sha256cu.m_pad_pars.block_512[15][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06288_));
 sky130_fd_sc_hd__a21oi_1 _12622_ (.A1(_01966_),
    .A2(_04938_),
    .B1(_06288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_2 _12623_ (.A(_06270_),
    .B(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06289_));
 sky130_fd_sc_hd__and2_1 _12624_ (.A(\sha256cu.m_pad_pars.block_512[16][0] ),
    .B(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _12625_ (.A(_06290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01065_));
 sky130_fd_sc_hd__and2_1 _12626_ (.A(\sha256cu.m_pad_pars.block_512[16][1] ),
    .B(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06291_));
 sky130_fd_sc_hd__clkbuf_1 _12627_ (.A(_06291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01066_));
 sky130_fd_sc_hd__and2_1 _12628_ (.A(\sha256cu.m_pad_pars.block_512[16][2] ),
    .B(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06292_));
 sky130_fd_sc_hd__clkbuf_1 _12629_ (.A(_06292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01067_));
 sky130_fd_sc_hd__and2_1 _12630_ (.A(\sha256cu.m_pad_pars.block_512[16][3] ),
    .B(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06293_));
 sky130_fd_sc_hd__clkbuf_1 _12631_ (.A(_06293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01068_));
 sky130_fd_sc_hd__and2_1 _12632_ (.A(\sha256cu.m_pad_pars.block_512[16][4] ),
    .B(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06294_));
 sky130_fd_sc_hd__clkbuf_1 _12633_ (.A(_06294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01069_));
 sky130_fd_sc_hd__and2_1 _12634_ (.A(\sha256cu.m_pad_pars.block_512[16][5] ),
    .B(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06295_));
 sky130_fd_sc_hd__clkbuf_1 _12635_ (.A(_06295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01070_));
 sky130_fd_sc_hd__and2_1 _12636_ (.A(\sha256cu.m_pad_pars.block_512[16][6] ),
    .B(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06296_));
 sky130_fd_sc_hd__clkbuf_1 _12637_ (.A(_06296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _12638_ (.A0(\sha256cu.m_pad_pars.block_512[16][7] ),
    .A1(_05413_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06297_));
 sky130_fd_sc_hd__clkbuf_1 _12639_ (.A(_06297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01072_));
 sky130_fd_sc_hd__or2_2 _12640_ (.A(_01912_),
    .B(_05137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06298_));
 sky130_fd_sc_hd__and2_1 _12641_ (.A(\sha256cu.m_pad_pars.block_512[17][0] ),
    .B(_06298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06299_));
 sky130_fd_sc_hd__clkbuf_1 _12642_ (.A(_06299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01073_));
 sky130_fd_sc_hd__and2_1 _12643_ (.A(\sha256cu.m_pad_pars.block_512[17][1] ),
    .B(_06298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06300_));
 sky130_fd_sc_hd__clkbuf_1 _12644_ (.A(_06300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01074_));
 sky130_fd_sc_hd__and2_1 _12645_ (.A(\sha256cu.m_pad_pars.block_512[17][2] ),
    .B(_06298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06301_));
 sky130_fd_sc_hd__clkbuf_1 _12646_ (.A(_06301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01075_));
 sky130_fd_sc_hd__and2_1 _12647_ (.A(\sha256cu.m_pad_pars.block_512[17][3] ),
    .B(_06298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06302_));
 sky130_fd_sc_hd__clkbuf_1 _12648_ (.A(_06302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01076_));
 sky130_fd_sc_hd__and2_1 _12649_ (.A(\sha256cu.m_pad_pars.block_512[17][4] ),
    .B(_06298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06303_));
 sky130_fd_sc_hd__clkbuf_1 _12650_ (.A(_06303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01077_));
 sky130_fd_sc_hd__and2_1 _12651_ (.A(\sha256cu.m_pad_pars.block_512[17][5] ),
    .B(_06298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06304_));
 sky130_fd_sc_hd__clkbuf_1 _12652_ (.A(_06304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01078_));
 sky130_fd_sc_hd__and2_1 _12653_ (.A(\sha256cu.m_pad_pars.block_512[17][6] ),
    .B(_06298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06305_));
 sky130_fd_sc_hd__clkbuf_1 _12654_ (.A(_06305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _12655_ (.A0(\sha256cu.m_pad_pars.block_512[17][7] ),
    .A1(_05266_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06306_));
 sky130_fd_sc_hd__clkbuf_1 _12656_ (.A(_06306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01080_));
 sky130_fd_sc_hd__or3_4 _12657_ (.A(_06251_),
    .B(_05081_),
    .C(_04994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06307_));
 sky130_fd_sc_hd__and2_1 _12658_ (.A(\sha256cu.m_pad_pars.block_512[18][0] ),
    .B(_06307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06308_));
 sky130_fd_sc_hd__clkbuf_1 _12659_ (.A(_06308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01081_));
 sky130_fd_sc_hd__and2_1 _12660_ (.A(\sha256cu.m_pad_pars.block_512[18][1] ),
    .B(_06307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06309_));
 sky130_fd_sc_hd__clkbuf_1 _12661_ (.A(_06309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01082_));
 sky130_fd_sc_hd__and2_1 _12662_ (.A(\sha256cu.m_pad_pars.block_512[18][2] ),
    .B(_06307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06310_));
 sky130_fd_sc_hd__clkbuf_1 _12663_ (.A(_06310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01083_));
 sky130_fd_sc_hd__and2_1 _12664_ (.A(\sha256cu.m_pad_pars.block_512[18][3] ),
    .B(_06307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06311_));
 sky130_fd_sc_hd__clkbuf_1 _12665_ (.A(_06311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01084_));
 sky130_fd_sc_hd__and2_1 _12666_ (.A(\sha256cu.m_pad_pars.block_512[18][4] ),
    .B(_06307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06312_));
 sky130_fd_sc_hd__clkbuf_1 _12667_ (.A(_06312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01085_));
 sky130_fd_sc_hd__and2_1 _12668_ (.A(\sha256cu.m_pad_pars.block_512[18][5] ),
    .B(_06307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06313_));
 sky130_fd_sc_hd__clkbuf_1 _12669_ (.A(_06313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01086_));
 sky130_fd_sc_hd__and2_1 _12670_ (.A(\sha256cu.m_pad_pars.block_512[18][6] ),
    .B(_06307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06314_));
 sky130_fd_sc_hd__clkbuf_1 _12671_ (.A(_06314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _12672_ (.A0(\sha256cu.m_pad_pars.block_512[18][7] ),
    .A1(_05108_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_1 _12673_ (.A(_06315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01088_));
 sky130_fd_sc_hd__or2_2 _12674_ (.A(_01912_),
    .B(_04830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06316_));
 sky130_fd_sc_hd__and2_1 _12675_ (.A(\sha256cu.m_pad_pars.block_512[19][0] ),
    .B(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06317_));
 sky130_fd_sc_hd__clkbuf_1 _12676_ (.A(_06317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01089_));
 sky130_fd_sc_hd__and2_1 _12677_ (.A(\sha256cu.m_pad_pars.block_512[19][1] ),
    .B(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06318_));
 sky130_fd_sc_hd__clkbuf_1 _12678_ (.A(_06318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01090_));
 sky130_fd_sc_hd__and2_1 _12679_ (.A(\sha256cu.m_pad_pars.block_512[19][2] ),
    .B(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06319_));
 sky130_fd_sc_hd__clkbuf_1 _12680_ (.A(_06319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01091_));
 sky130_fd_sc_hd__and2_1 _12681_ (.A(\sha256cu.m_pad_pars.block_512[19][3] ),
    .B(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06320_));
 sky130_fd_sc_hd__clkbuf_1 _12682_ (.A(_06320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01092_));
 sky130_fd_sc_hd__and2_1 _12683_ (.A(\sha256cu.m_pad_pars.block_512[19][4] ),
    .B(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_1 _12684_ (.A(_06321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01093_));
 sky130_fd_sc_hd__and2_1 _12685_ (.A(\sha256cu.m_pad_pars.block_512[19][5] ),
    .B(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06322_));
 sky130_fd_sc_hd__clkbuf_1 _12686_ (.A(_06322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01094_));
 sky130_fd_sc_hd__and2_1 _12687_ (.A(\sha256cu.m_pad_pars.block_512[19][6] ),
    .B(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06323_));
 sky130_fd_sc_hd__clkbuf_1 _12688_ (.A(_06323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(\sha256cu.m_pad_pars.block_512[19][7] ),
    .A1(_04943_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06324_));
 sky130_fd_sc_hd__clkbuf_1 _12690_ (.A(_06324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01096_));
 sky130_fd_sc_hd__or3_4 _12691_ (.A(_06251_),
    .B(_05081_),
    .C(_05292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06325_));
 sky130_fd_sc_hd__and2_1 _12692_ (.A(\sha256cu.m_pad_pars.block_512[20][0] ),
    .B(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_1 _12693_ (.A(_06326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01097_));
 sky130_fd_sc_hd__and2_1 _12694_ (.A(\sha256cu.m_pad_pars.block_512[20][1] ),
    .B(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06327_));
 sky130_fd_sc_hd__clkbuf_1 _12695_ (.A(_06327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01098_));
 sky130_fd_sc_hd__and2_1 _12696_ (.A(\sha256cu.m_pad_pars.block_512[20][2] ),
    .B(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06328_));
 sky130_fd_sc_hd__clkbuf_1 _12697_ (.A(_06328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01099_));
 sky130_fd_sc_hd__and2_1 _12698_ (.A(\sha256cu.m_pad_pars.block_512[20][3] ),
    .B(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06329_));
 sky130_fd_sc_hd__clkbuf_1 _12699_ (.A(_06329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01100_));
 sky130_fd_sc_hd__and2_1 _12700_ (.A(\sha256cu.m_pad_pars.block_512[20][4] ),
    .B(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06330_));
 sky130_fd_sc_hd__clkbuf_1 _12701_ (.A(_06330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01101_));
 sky130_fd_sc_hd__and2_1 _12702_ (.A(\sha256cu.m_pad_pars.block_512[20][5] ),
    .B(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06331_));
 sky130_fd_sc_hd__clkbuf_1 _12703_ (.A(_06331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01102_));
 sky130_fd_sc_hd__and2_1 _12704_ (.A(\sha256cu.m_pad_pars.block_512[20][6] ),
    .B(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06332_));
 sky130_fd_sc_hd__clkbuf_1 _12705_ (.A(_06332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _12706_ (.A0(\sha256cu.m_pad_pars.block_512[20][7] ),
    .A1(_05396_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06333_));
 sky130_fd_sc_hd__clkbuf_1 _12707_ (.A(_06333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01104_));
 sky130_fd_sc_hd__nand2_2 _12708_ (.A(_06270_),
    .B(_05156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06334_));
 sky130_fd_sc_hd__and2_1 _12709_ (.A(\sha256cu.m_pad_pars.block_512[21][0] ),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06335_));
 sky130_fd_sc_hd__clkbuf_1 _12710_ (.A(_06335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01105_));
 sky130_fd_sc_hd__and2_1 _12711_ (.A(\sha256cu.m_pad_pars.block_512[21][1] ),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06336_));
 sky130_fd_sc_hd__clkbuf_1 _12712_ (.A(_06336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01106_));
 sky130_fd_sc_hd__and2_1 _12713_ (.A(\sha256cu.m_pad_pars.block_512[21][2] ),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06337_));
 sky130_fd_sc_hd__clkbuf_1 _12714_ (.A(_06337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01107_));
 sky130_fd_sc_hd__and2_1 _12715_ (.A(\sha256cu.m_pad_pars.block_512[21][3] ),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06338_));
 sky130_fd_sc_hd__clkbuf_1 _12716_ (.A(_06338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01108_));
 sky130_fd_sc_hd__and2_1 _12717_ (.A(\sha256cu.m_pad_pars.block_512[21][4] ),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06339_));
 sky130_fd_sc_hd__clkbuf_1 _12718_ (.A(_06339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01109_));
 sky130_fd_sc_hd__and2_1 _12719_ (.A(\sha256cu.m_pad_pars.block_512[21][5] ),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06340_));
 sky130_fd_sc_hd__clkbuf_1 _12720_ (.A(_06340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01110_));
 sky130_fd_sc_hd__and2_1 _12721_ (.A(\sha256cu.m_pad_pars.block_512[21][6] ),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06341_));
 sky130_fd_sc_hd__clkbuf_1 _12722_ (.A(_06341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _12723_ (.A0(\sha256cu.m_pad_pars.block_512[21][7] ),
    .A1(_05236_),
    .S(_06249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06342_));
 sky130_fd_sc_hd__clkbuf_1 _12724_ (.A(_06342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01112_));
 sky130_fd_sc_hd__o21ai_4 _12725_ (.A1(_05011_),
    .A2(_05012_),
    .B1(_06270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06343_));
 sky130_fd_sc_hd__and2_1 _12726_ (.A(\sha256cu.m_pad_pars.block_512[22][0] ),
    .B(_06343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06344_));
 sky130_fd_sc_hd__clkbuf_1 _12727_ (.A(_06344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01113_));
 sky130_fd_sc_hd__and2_1 _12728_ (.A(\sha256cu.m_pad_pars.block_512[22][1] ),
    .B(_06343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06345_));
 sky130_fd_sc_hd__clkbuf_1 _12729_ (.A(_06345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01114_));
 sky130_fd_sc_hd__and2_1 _12730_ (.A(\sha256cu.m_pad_pars.block_512[22][2] ),
    .B(_06343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06346_));
 sky130_fd_sc_hd__clkbuf_1 _12731_ (.A(_06346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01115_));
 sky130_fd_sc_hd__and2_1 _12732_ (.A(\sha256cu.m_pad_pars.block_512[22][3] ),
    .B(_06343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06347_));
 sky130_fd_sc_hd__clkbuf_1 _12733_ (.A(_06347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01116_));
 sky130_fd_sc_hd__and2_1 _12734_ (.A(\sha256cu.m_pad_pars.block_512[22][4] ),
    .B(_06343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06348_));
 sky130_fd_sc_hd__clkbuf_1 _12735_ (.A(_06348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01117_));
 sky130_fd_sc_hd__and2_1 _12736_ (.A(\sha256cu.m_pad_pars.block_512[22][5] ),
    .B(_06343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06349_));
 sky130_fd_sc_hd__clkbuf_1 _12737_ (.A(_06349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01118_));
 sky130_fd_sc_hd__and2_1 _12738_ (.A(\sha256cu.m_pad_pars.block_512[22][6] ),
    .B(_06343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_1 _12739_ (.A(_06350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01119_));
 sky130_fd_sc_hd__buf_4 _12740_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06351_));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(\sha256cu.m_pad_pars.block_512[22][7] ),
    .A1(_05111_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06352_));
 sky130_fd_sc_hd__clkbuf_1 _12742_ (.A(_06352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01120_));
 sky130_fd_sc_hd__or2_2 _12743_ (.A(_01912_),
    .B(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06353_));
 sky130_fd_sc_hd__and2_1 _12744_ (.A(\sha256cu.m_pad_pars.block_512[23][0] ),
    .B(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_1 _12745_ (.A(_06354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01121_));
 sky130_fd_sc_hd__and2_1 _12746_ (.A(\sha256cu.m_pad_pars.block_512[23][1] ),
    .B(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06355_));
 sky130_fd_sc_hd__clkbuf_1 _12747_ (.A(_06355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01122_));
 sky130_fd_sc_hd__and2_1 _12748_ (.A(\sha256cu.m_pad_pars.block_512[23][2] ),
    .B(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _12749_ (.A(_06356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01123_));
 sky130_fd_sc_hd__and2_1 _12750_ (.A(\sha256cu.m_pad_pars.block_512[23][3] ),
    .B(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06357_));
 sky130_fd_sc_hd__clkbuf_1 _12751_ (.A(_06357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01124_));
 sky130_fd_sc_hd__and2_1 _12752_ (.A(\sha256cu.m_pad_pars.block_512[23][4] ),
    .B(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06358_));
 sky130_fd_sc_hd__clkbuf_1 _12753_ (.A(_06358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01125_));
 sky130_fd_sc_hd__and2_1 _12754_ (.A(\sha256cu.m_pad_pars.block_512[23][5] ),
    .B(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06359_));
 sky130_fd_sc_hd__clkbuf_1 _12755_ (.A(_06359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01126_));
 sky130_fd_sc_hd__and2_1 _12756_ (.A(\sha256cu.m_pad_pars.block_512[23][6] ),
    .B(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06360_));
 sky130_fd_sc_hd__clkbuf_1 _12757_ (.A(_06360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _12758_ (.A0(\sha256cu.m_pad_pars.block_512[23][7] ),
    .A1(_04927_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06361_));
 sky130_fd_sc_hd__clkbuf_1 _12759_ (.A(_06361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01128_));
 sky130_fd_sc_hd__or3_4 _12760_ (.A(_06251_),
    .B(_05081_),
    .C(_05276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06362_));
 sky130_fd_sc_hd__and2_1 _12761_ (.A(\sha256cu.m_pad_pars.block_512[24][0] ),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06363_));
 sky130_fd_sc_hd__clkbuf_1 _12762_ (.A(_06363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01129_));
 sky130_fd_sc_hd__and2_1 _12763_ (.A(\sha256cu.m_pad_pars.block_512[24][1] ),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_1 _12764_ (.A(_06364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01130_));
 sky130_fd_sc_hd__and2_1 _12765_ (.A(\sha256cu.m_pad_pars.block_512[24][2] ),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06365_));
 sky130_fd_sc_hd__clkbuf_1 _12766_ (.A(_06365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01131_));
 sky130_fd_sc_hd__and2_1 _12767_ (.A(\sha256cu.m_pad_pars.block_512[24][3] ),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _12768_ (.A(_06366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01132_));
 sky130_fd_sc_hd__and2_1 _12769_ (.A(\sha256cu.m_pad_pars.block_512[24][4] ),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06367_));
 sky130_fd_sc_hd__clkbuf_1 _12770_ (.A(_06367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01133_));
 sky130_fd_sc_hd__and2_1 _12771_ (.A(\sha256cu.m_pad_pars.block_512[24][5] ),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06368_));
 sky130_fd_sc_hd__clkbuf_1 _12772_ (.A(_06368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01134_));
 sky130_fd_sc_hd__and2_1 _12773_ (.A(\sha256cu.m_pad_pars.block_512[24][6] ),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06369_));
 sky130_fd_sc_hd__clkbuf_1 _12774_ (.A(_06369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _12775_ (.A0(\sha256cu.m_pad_pars.block_512[24][7] ),
    .A1(_05405_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06370_));
 sky130_fd_sc_hd__clkbuf_1 _12776_ (.A(_06370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01136_));
 sky130_fd_sc_hd__or3_2 _12777_ (.A(_06251_),
    .B(_05081_),
    .C(_05130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06371_));
 sky130_fd_sc_hd__and2_1 _12778_ (.A(\sha256cu.m_pad_pars.block_512[25][0] ),
    .B(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _12779_ (.A(_06372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01137_));
 sky130_fd_sc_hd__and2_1 _12780_ (.A(\sha256cu.m_pad_pars.block_512[25][1] ),
    .B(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06373_));
 sky130_fd_sc_hd__clkbuf_1 _12781_ (.A(_06373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01138_));
 sky130_fd_sc_hd__and2_1 _12782_ (.A(\sha256cu.m_pad_pars.block_512[25][2] ),
    .B(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_1 _12783_ (.A(_06374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01139_));
 sky130_fd_sc_hd__and2_1 _12784_ (.A(\sha256cu.m_pad_pars.block_512[25][3] ),
    .B(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06375_));
 sky130_fd_sc_hd__clkbuf_1 _12785_ (.A(_06375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01140_));
 sky130_fd_sc_hd__and2_1 _12786_ (.A(\sha256cu.m_pad_pars.block_512[25][4] ),
    .B(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06376_));
 sky130_fd_sc_hd__clkbuf_1 _12787_ (.A(_06376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01141_));
 sky130_fd_sc_hd__and2_1 _12788_ (.A(\sha256cu.m_pad_pars.block_512[25][5] ),
    .B(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_1 _12789_ (.A(_06377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01142_));
 sky130_fd_sc_hd__and2_1 _12790_ (.A(\sha256cu.m_pad_pars.block_512[25][6] ),
    .B(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _12791_ (.A(_06378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _12792_ (.A0(\sha256cu.m_pad_pars.block_512[25][7] ),
    .A1(_05243_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06379_));
 sky130_fd_sc_hd__clkbuf_1 _12793_ (.A(_06379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01144_));
 sky130_fd_sc_hd__or3_2 _12794_ (.A(_06251_),
    .B(_05081_),
    .C(_04961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06380_));
 sky130_fd_sc_hd__and2_1 _12795_ (.A(\sha256cu.m_pad_pars.block_512[26][0] ),
    .B(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06381_));
 sky130_fd_sc_hd__clkbuf_1 _12796_ (.A(_06381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01145_));
 sky130_fd_sc_hd__and2_1 _12797_ (.A(\sha256cu.m_pad_pars.block_512[26][1] ),
    .B(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06382_));
 sky130_fd_sc_hd__clkbuf_1 _12798_ (.A(_06382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01146_));
 sky130_fd_sc_hd__and2_1 _12799_ (.A(\sha256cu.m_pad_pars.block_512[26][2] ),
    .B(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06383_));
 sky130_fd_sc_hd__clkbuf_1 _12800_ (.A(_06383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01147_));
 sky130_fd_sc_hd__and2_1 _12801_ (.A(\sha256cu.m_pad_pars.block_512[26][3] ),
    .B(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06384_));
 sky130_fd_sc_hd__clkbuf_1 _12802_ (.A(_06384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01148_));
 sky130_fd_sc_hd__and2_1 _12803_ (.A(\sha256cu.m_pad_pars.block_512[26][4] ),
    .B(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06385_));
 sky130_fd_sc_hd__clkbuf_1 _12804_ (.A(_06385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01149_));
 sky130_fd_sc_hd__and2_1 _12805_ (.A(\sha256cu.m_pad_pars.block_512[26][5] ),
    .B(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06386_));
 sky130_fd_sc_hd__clkbuf_1 _12806_ (.A(_06386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01150_));
 sky130_fd_sc_hd__and2_1 _12807_ (.A(\sha256cu.m_pad_pars.block_512[26][6] ),
    .B(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06387_));
 sky130_fd_sc_hd__clkbuf_1 _12808_ (.A(_06387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(\sha256cu.m_pad_pars.block_512[26][7] ),
    .A1(_05083_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_1 _12810_ (.A(_06388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01152_));
 sky130_fd_sc_hd__or3_4 _12811_ (.A(_06251_),
    .B(_05081_),
    .C(_04754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06389_));
 sky130_fd_sc_hd__and2_1 _12812_ (.A(\sha256cu.m_pad_pars.block_512[27][0] ),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06390_));
 sky130_fd_sc_hd__clkbuf_1 _12813_ (.A(_06390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01153_));
 sky130_fd_sc_hd__and2_1 _12814_ (.A(\sha256cu.m_pad_pars.block_512[27][1] ),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06391_));
 sky130_fd_sc_hd__clkbuf_1 _12815_ (.A(_06391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01154_));
 sky130_fd_sc_hd__and2_1 _12816_ (.A(\sha256cu.m_pad_pars.block_512[27][2] ),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_1 _12817_ (.A(_06392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01155_));
 sky130_fd_sc_hd__and2_1 _12818_ (.A(\sha256cu.m_pad_pars.block_512[27][3] ),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06393_));
 sky130_fd_sc_hd__clkbuf_1 _12819_ (.A(_06393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01156_));
 sky130_fd_sc_hd__and2_1 _12820_ (.A(\sha256cu.m_pad_pars.block_512[27][4] ),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_1 _12821_ (.A(_06394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01157_));
 sky130_fd_sc_hd__and2_1 _12822_ (.A(\sha256cu.m_pad_pars.block_512[27][5] ),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06395_));
 sky130_fd_sc_hd__clkbuf_1 _12823_ (.A(_06395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01158_));
 sky130_fd_sc_hd__and2_1 _12824_ (.A(\sha256cu.m_pad_pars.block_512[27][6] ),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06396_));
 sky130_fd_sc_hd__clkbuf_1 _12825_ (.A(_06396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _12826_ (.A0(\sha256cu.m_pad_pars.block_512[27][7] ),
    .A1(_04945_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_1 _12827_ (.A(_06397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01160_));
 sky130_fd_sc_hd__or3_2 _12828_ (.A(_06251_),
    .B(_05081_),
    .C(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06398_));
 sky130_fd_sc_hd__and2_1 _12829_ (.A(\sha256cu.m_pad_pars.block_512[28][0] ),
    .B(_06398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06399_));
 sky130_fd_sc_hd__clkbuf_1 _12830_ (.A(_06399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01161_));
 sky130_fd_sc_hd__and2_1 _12831_ (.A(\sha256cu.m_pad_pars.block_512[28][1] ),
    .B(_06398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_1 _12832_ (.A(_06400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01162_));
 sky130_fd_sc_hd__and2_1 _12833_ (.A(\sha256cu.m_pad_pars.block_512[28][2] ),
    .B(_06398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06401_));
 sky130_fd_sc_hd__clkbuf_1 _12834_ (.A(_06401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01163_));
 sky130_fd_sc_hd__and2_1 _12835_ (.A(\sha256cu.m_pad_pars.block_512[28][3] ),
    .B(_06398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06402_));
 sky130_fd_sc_hd__clkbuf_1 _12836_ (.A(_06402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01164_));
 sky130_fd_sc_hd__and2_1 _12837_ (.A(\sha256cu.m_pad_pars.block_512[28][4] ),
    .B(_06398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_1 _12838_ (.A(_06403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01165_));
 sky130_fd_sc_hd__and2_1 _12839_ (.A(\sha256cu.m_pad_pars.block_512[28][5] ),
    .B(_06398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06404_));
 sky130_fd_sc_hd__clkbuf_1 _12840_ (.A(_06404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01166_));
 sky130_fd_sc_hd__and2_1 _12841_ (.A(\sha256cu.m_pad_pars.block_512[28][6] ),
    .B(_06398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06405_));
 sky130_fd_sc_hd__clkbuf_1 _12842_ (.A(_06405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(\sha256cu.m_pad_pars.block_512[28][7] ),
    .A1(_05388_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_1 _12844_ (.A(_06406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01168_));
 sky130_fd_sc_hd__or3_4 _12845_ (.A(_06251_),
    .B(_05081_),
    .C(_05124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06407_));
 sky130_fd_sc_hd__and2_1 _12846_ (.A(\sha256cu.m_pad_pars.block_512[29][0] ),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06408_));
 sky130_fd_sc_hd__clkbuf_1 _12847_ (.A(_06408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01169_));
 sky130_fd_sc_hd__and2_1 _12848_ (.A(\sha256cu.m_pad_pars.block_512[29][1] ),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06409_));
 sky130_fd_sc_hd__clkbuf_1 _12849_ (.A(_06409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01170_));
 sky130_fd_sc_hd__and2_1 _12850_ (.A(\sha256cu.m_pad_pars.block_512[29][2] ),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06410_));
 sky130_fd_sc_hd__clkbuf_1 _12851_ (.A(_06410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01171_));
 sky130_fd_sc_hd__and2_1 _12852_ (.A(\sha256cu.m_pad_pars.block_512[29][3] ),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06411_));
 sky130_fd_sc_hd__clkbuf_1 _12853_ (.A(_06411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01172_));
 sky130_fd_sc_hd__and2_1 _12854_ (.A(\sha256cu.m_pad_pars.block_512[29][4] ),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_1 _12855_ (.A(_06412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01173_));
 sky130_fd_sc_hd__and2_1 _12856_ (.A(\sha256cu.m_pad_pars.block_512[29][5] ),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06413_));
 sky130_fd_sc_hd__clkbuf_1 _12857_ (.A(_06413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01174_));
 sky130_fd_sc_hd__and2_1 _12858_ (.A(\sha256cu.m_pad_pars.block_512[29][6] ),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06414_));
 sky130_fd_sc_hd__clkbuf_1 _12859_ (.A(_06414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(\sha256cu.m_pad_pars.block_512[29][7] ),
    .A1(_05250_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_1 _12861_ (.A(_06415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01176_));
 sky130_fd_sc_hd__or3_2 _12862_ (.A(_02111_),
    .B(_05081_),
    .C(_04975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06416_));
 sky130_fd_sc_hd__and2_1 _12863_ (.A(\sha256cu.m_pad_pars.block_512[30][0] ),
    .B(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06417_));
 sky130_fd_sc_hd__clkbuf_1 _12864_ (.A(_06417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01177_));
 sky130_fd_sc_hd__and2_1 _12865_ (.A(\sha256cu.m_pad_pars.block_512[30][1] ),
    .B(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06418_));
 sky130_fd_sc_hd__clkbuf_1 _12866_ (.A(_06418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01178_));
 sky130_fd_sc_hd__and2_1 _12867_ (.A(\sha256cu.m_pad_pars.block_512[30][2] ),
    .B(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06419_));
 sky130_fd_sc_hd__clkbuf_1 _12868_ (.A(_06419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01179_));
 sky130_fd_sc_hd__and2_1 _12869_ (.A(\sha256cu.m_pad_pars.block_512[30][3] ),
    .B(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06420_));
 sky130_fd_sc_hd__clkbuf_1 _12870_ (.A(_06420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01180_));
 sky130_fd_sc_hd__and2_1 _12871_ (.A(\sha256cu.m_pad_pars.block_512[30][4] ),
    .B(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06421_));
 sky130_fd_sc_hd__clkbuf_1 _12872_ (.A(_06421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01181_));
 sky130_fd_sc_hd__and2_1 _12873_ (.A(\sha256cu.m_pad_pars.block_512[30][5] ),
    .B(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06422_));
 sky130_fd_sc_hd__clkbuf_1 _12874_ (.A(_06422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01182_));
 sky130_fd_sc_hd__and2_1 _12875_ (.A(\sha256cu.m_pad_pars.block_512[30][6] ),
    .B(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06423_));
 sky130_fd_sc_hd__clkbuf_1 _12876_ (.A(_06423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _12877_ (.A0(\sha256cu.m_pad_pars.block_512[30][7] ),
    .A1(_05102_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06424_));
 sky130_fd_sc_hd__clkbuf_1 _12878_ (.A(_06424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01184_));
 sky130_fd_sc_hd__or3_2 _12879_ (.A(_02111_),
    .B(_04705_),
    .C(_04809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06425_));
 sky130_fd_sc_hd__and2_1 _12880_ (.A(\sha256cu.m_pad_pars.block_512[31][0] ),
    .B(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_1 _12881_ (.A(_06426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01185_));
 sky130_fd_sc_hd__and2_1 _12882_ (.A(\sha256cu.m_pad_pars.block_512[31][1] ),
    .B(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06427_));
 sky130_fd_sc_hd__clkbuf_1 _12883_ (.A(_06427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01186_));
 sky130_fd_sc_hd__and2_1 _12884_ (.A(\sha256cu.m_pad_pars.block_512[31][2] ),
    .B(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06428_));
 sky130_fd_sc_hd__clkbuf_1 _12885_ (.A(_06428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01187_));
 sky130_fd_sc_hd__and2_1 _12886_ (.A(\sha256cu.m_pad_pars.block_512[31][3] ),
    .B(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06429_));
 sky130_fd_sc_hd__clkbuf_1 _12887_ (.A(_06429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01188_));
 sky130_fd_sc_hd__and2_1 _12888_ (.A(\sha256cu.m_pad_pars.block_512[31][4] ),
    .B(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_1 _12889_ (.A(_06430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01189_));
 sky130_fd_sc_hd__and2_1 _12890_ (.A(\sha256cu.m_pad_pars.block_512[31][5] ),
    .B(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06431_));
 sky130_fd_sc_hd__clkbuf_1 _12891_ (.A(_06431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01190_));
 sky130_fd_sc_hd__and2_1 _12892_ (.A(\sha256cu.m_pad_pars.block_512[31][6] ),
    .B(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06432_));
 sky130_fd_sc_hd__clkbuf_1 _12893_ (.A(_06432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(\sha256cu.m_pad_pars.block_512[31][7] ),
    .A1(_04911_),
    .S(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06433_));
 sky130_fd_sc_hd__clkbuf_1 _12895_ (.A(_06433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01192_));
 sky130_fd_sc_hd__or2_2 _12896_ (.A(_01912_),
    .B(_05305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06434_));
 sky130_fd_sc_hd__and2_1 _12897_ (.A(\sha256cu.m_pad_pars.block_512[32][0] ),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06435_));
 sky130_fd_sc_hd__clkbuf_1 _12898_ (.A(_06435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01193_));
 sky130_fd_sc_hd__and2_1 _12899_ (.A(\sha256cu.m_pad_pars.block_512[32][1] ),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06436_));
 sky130_fd_sc_hd__clkbuf_1 _12900_ (.A(_06436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01194_));
 sky130_fd_sc_hd__and2_1 _12901_ (.A(\sha256cu.m_pad_pars.block_512[32][2] ),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06437_));
 sky130_fd_sc_hd__clkbuf_1 _12902_ (.A(_06437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01195_));
 sky130_fd_sc_hd__and2_1 _12903_ (.A(\sha256cu.m_pad_pars.block_512[32][3] ),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06438_));
 sky130_fd_sc_hd__clkbuf_1 _12904_ (.A(_06438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01196_));
 sky130_fd_sc_hd__and2_1 _12905_ (.A(\sha256cu.m_pad_pars.block_512[32][4] ),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_1 _12906_ (.A(_06439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01197_));
 sky130_fd_sc_hd__and2_1 _12907_ (.A(\sha256cu.m_pad_pars.block_512[32][5] ),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06440_));
 sky130_fd_sc_hd__clkbuf_1 _12908_ (.A(_06440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01198_));
 sky130_fd_sc_hd__and2_1 _12909_ (.A(\sha256cu.m_pad_pars.block_512[32][6] ),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06441_));
 sky130_fd_sc_hd__clkbuf_1 _12910_ (.A(_06441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01199_));
 sky130_fd_sc_hd__buf_4 _12911_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06442_));
 sky130_fd_sc_hd__mux2_1 _12912_ (.A0(\sha256cu.m_pad_pars.block_512[32][7] ),
    .A1(_05394_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06443_));
 sky130_fd_sc_hd__clkbuf_1 _12913_ (.A(_06443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01200_));
 sky130_fd_sc_hd__or2_2 _12914_ (.A(_01912_),
    .B(_05146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06444_));
 sky130_fd_sc_hd__and2_1 _12915_ (.A(\sha256cu.m_pad_pars.block_512[33][0] ),
    .B(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06445_));
 sky130_fd_sc_hd__clkbuf_1 _12916_ (.A(_06445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01201_));
 sky130_fd_sc_hd__and2_1 _12917_ (.A(\sha256cu.m_pad_pars.block_512[33][1] ),
    .B(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06446_));
 sky130_fd_sc_hd__clkbuf_1 _12918_ (.A(_06446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01202_));
 sky130_fd_sc_hd__and2_1 _12919_ (.A(\sha256cu.m_pad_pars.block_512[33][2] ),
    .B(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06447_));
 sky130_fd_sc_hd__clkbuf_1 _12920_ (.A(_06447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01203_));
 sky130_fd_sc_hd__and2_1 _12921_ (.A(\sha256cu.m_pad_pars.block_512[33][3] ),
    .B(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06448_));
 sky130_fd_sc_hd__clkbuf_1 _12922_ (.A(_06448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01204_));
 sky130_fd_sc_hd__and2_1 _12923_ (.A(\sha256cu.m_pad_pars.block_512[33][4] ),
    .B(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06449_));
 sky130_fd_sc_hd__clkbuf_1 _12924_ (.A(_06449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01205_));
 sky130_fd_sc_hd__and2_1 _12925_ (.A(\sha256cu.m_pad_pars.block_512[33][5] ),
    .B(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06450_));
 sky130_fd_sc_hd__clkbuf_1 _12926_ (.A(_06450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01206_));
 sky130_fd_sc_hd__and2_1 _12927_ (.A(\sha256cu.m_pad_pars.block_512[33][6] ),
    .B(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06451_));
 sky130_fd_sc_hd__clkbuf_1 _12928_ (.A(_06451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _12929_ (.A0(\sha256cu.m_pad_pars.block_512[33][7] ),
    .A1(_05267_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06452_));
 sky130_fd_sc_hd__clkbuf_1 _12930_ (.A(_06452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01208_));
 sky130_fd_sc_hd__nand2_2 _12931_ (.A(_06270_),
    .B(_04995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06453_));
 sky130_fd_sc_hd__and2_1 _12932_ (.A(\sha256cu.m_pad_pars.block_512[34][0] ),
    .B(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06454_));
 sky130_fd_sc_hd__clkbuf_1 _12933_ (.A(_06454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01209_));
 sky130_fd_sc_hd__and2_1 _12934_ (.A(\sha256cu.m_pad_pars.block_512[34][1] ),
    .B(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06455_));
 sky130_fd_sc_hd__clkbuf_1 _12935_ (.A(_06455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01210_));
 sky130_fd_sc_hd__and2_1 _12936_ (.A(\sha256cu.m_pad_pars.block_512[34][2] ),
    .B(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06456_));
 sky130_fd_sc_hd__clkbuf_1 _12937_ (.A(_06456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01211_));
 sky130_fd_sc_hd__and2_1 _12938_ (.A(\sha256cu.m_pad_pars.block_512[34][3] ),
    .B(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06457_));
 sky130_fd_sc_hd__clkbuf_1 _12939_ (.A(_06457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01212_));
 sky130_fd_sc_hd__and2_1 _12940_ (.A(\sha256cu.m_pad_pars.block_512[34][4] ),
    .B(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06458_));
 sky130_fd_sc_hd__clkbuf_1 _12941_ (.A(_06458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01213_));
 sky130_fd_sc_hd__and2_1 _12942_ (.A(\sha256cu.m_pad_pars.block_512[34][5] ),
    .B(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06459_));
 sky130_fd_sc_hd__clkbuf_1 _12943_ (.A(_06459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01214_));
 sky130_fd_sc_hd__and2_1 _12944_ (.A(\sha256cu.m_pad_pars.block_512[34][6] ),
    .B(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_1 _12945_ (.A(_06460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01215_));
 sky130_fd_sc_hd__nor2_1 _12946_ (.A(_03288_),
    .B(\sha256cu.m_pad_pars.block_512[34][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06461_));
 sky130_fd_sc_hd__a21oi_1 _12947_ (.A1(_01966_),
    .A2(_05121_),
    .B1(_06461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01216_));
 sky130_fd_sc_hd__nand2_2 _12948_ (.A(_06270_),
    .B(_04817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06462_));
 sky130_fd_sc_hd__and2_1 _12949_ (.A(\sha256cu.m_pad_pars.block_512[35][0] ),
    .B(_06462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06463_));
 sky130_fd_sc_hd__clkbuf_1 _12950_ (.A(_06463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01217_));
 sky130_fd_sc_hd__and2_1 _12951_ (.A(\sha256cu.m_pad_pars.block_512[35][1] ),
    .B(_06462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06464_));
 sky130_fd_sc_hd__clkbuf_1 _12952_ (.A(_06464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01218_));
 sky130_fd_sc_hd__and2_1 _12953_ (.A(\sha256cu.m_pad_pars.block_512[35][2] ),
    .B(_06462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06465_));
 sky130_fd_sc_hd__clkbuf_1 _12954_ (.A(_06465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01219_));
 sky130_fd_sc_hd__and2_1 _12955_ (.A(\sha256cu.m_pad_pars.block_512[35][3] ),
    .B(_06462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06466_));
 sky130_fd_sc_hd__clkbuf_1 _12956_ (.A(_06466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01220_));
 sky130_fd_sc_hd__and2_1 _12957_ (.A(\sha256cu.m_pad_pars.block_512[35][4] ),
    .B(_06462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06467_));
 sky130_fd_sc_hd__clkbuf_1 _12958_ (.A(_06467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01221_));
 sky130_fd_sc_hd__and2_1 _12959_ (.A(\sha256cu.m_pad_pars.block_512[35][5] ),
    .B(_06462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06468_));
 sky130_fd_sc_hd__clkbuf_1 _12960_ (.A(_06468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01222_));
 sky130_fd_sc_hd__and2_1 _12961_ (.A(\sha256cu.m_pad_pars.block_512[35][6] ),
    .B(_06462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06469_));
 sky130_fd_sc_hd__clkbuf_1 _12962_ (.A(_06469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _12963_ (.A0(\sha256cu.m_pad_pars.block_512[35][7] ),
    .A1(_04920_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06470_));
 sky130_fd_sc_hd__clkbuf_1 _12964_ (.A(_06470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01224_));
 sky130_fd_sc_hd__or2_2 _12965_ (.A(_01986_),
    .B(_05303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06471_));
 sky130_fd_sc_hd__and2_1 _12966_ (.A(\sha256cu.m_pad_pars.block_512[36][0] ),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06472_));
 sky130_fd_sc_hd__clkbuf_1 _12967_ (.A(_06472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01225_));
 sky130_fd_sc_hd__and2_1 _12968_ (.A(\sha256cu.m_pad_pars.block_512[36][1] ),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06473_));
 sky130_fd_sc_hd__clkbuf_1 _12969_ (.A(_06473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01226_));
 sky130_fd_sc_hd__and2_1 _12970_ (.A(\sha256cu.m_pad_pars.block_512[36][2] ),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06474_));
 sky130_fd_sc_hd__clkbuf_1 _12971_ (.A(_06474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01227_));
 sky130_fd_sc_hd__and2_1 _12972_ (.A(\sha256cu.m_pad_pars.block_512[36][3] ),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06475_));
 sky130_fd_sc_hd__clkbuf_1 _12973_ (.A(_06475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01228_));
 sky130_fd_sc_hd__and2_1 _12974_ (.A(\sha256cu.m_pad_pars.block_512[36][4] ),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06476_));
 sky130_fd_sc_hd__clkbuf_1 _12975_ (.A(_06476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01229_));
 sky130_fd_sc_hd__and2_1 _12976_ (.A(\sha256cu.m_pad_pars.block_512[36][5] ),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06477_));
 sky130_fd_sc_hd__clkbuf_1 _12977_ (.A(_06477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01230_));
 sky130_fd_sc_hd__and2_1 _12978_ (.A(\sha256cu.m_pad_pars.block_512[36][6] ),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06478_));
 sky130_fd_sc_hd__clkbuf_1 _12979_ (.A(_06478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _12980_ (.A0(\sha256cu.m_pad_pars.block_512[36][7] ),
    .A1(_05401_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06479_));
 sky130_fd_sc_hd__clkbuf_1 _12981_ (.A(_06479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01232_));
 sky130_fd_sc_hd__or3_2 _12982_ (.A(_02111_),
    .B(_04917_),
    .C(_05159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06480_));
 sky130_fd_sc_hd__and2_1 _12983_ (.A(\sha256cu.m_pad_pars.block_512[37][0] ),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06481_));
 sky130_fd_sc_hd__clkbuf_1 _12984_ (.A(_06481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01233_));
 sky130_fd_sc_hd__and2_1 _12985_ (.A(\sha256cu.m_pad_pars.block_512[37][1] ),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06482_));
 sky130_fd_sc_hd__clkbuf_1 _12986_ (.A(_06482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01234_));
 sky130_fd_sc_hd__and2_1 _12987_ (.A(\sha256cu.m_pad_pars.block_512[37][2] ),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06483_));
 sky130_fd_sc_hd__clkbuf_1 _12988_ (.A(_06483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01235_));
 sky130_fd_sc_hd__and2_1 _12989_ (.A(\sha256cu.m_pad_pars.block_512[37][3] ),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06484_));
 sky130_fd_sc_hd__clkbuf_1 _12990_ (.A(_06484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01236_));
 sky130_fd_sc_hd__and2_1 _12991_ (.A(\sha256cu.m_pad_pars.block_512[37][4] ),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06485_));
 sky130_fd_sc_hd__clkbuf_1 _12992_ (.A(_06485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01237_));
 sky130_fd_sc_hd__and2_1 _12993_ (.A(\sha256cu.m_pad_pars.block_512[37][5] ),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06486_));
 sky130_fd_sc_hd__clkbuf_1 _12994_ (.A(_06486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01238_));
 sky130_fd_sc_hd__and2_1 _12995_ (.A(\sha256cu.m_pad_pars.block_512[37][6] ),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06487_));
 sky130_fd_sc_hd__clkbuf_1 _12996_ (.A(_06487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _12997_ (.A0(\sha256cu.m_pad_pars.block_512[37][7] ),
    .A1(_05247_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06488_));
 sky130_fd_sc_hd__clkbuf_1 _12998_ (.A(_06488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01240_));
 sky130_fd_sc_hd__nand2_2 _12999_ (.A(_06270_),
    .B(_04971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06489_));
 sky130_fd_sc_hd__and2_1 _13000_ (.A(\sha256cu.m_pad_pars.block_512[38][0] ),
    .B(_06489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06490_));
 sky130_fd_sc_hd__clkbuf_1 _13001_ (.A(_06490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01241_));
 sky130_fd_sc_hd__and2_1 _13002_ (.A(\sha256cu.m_pad_pars.block_512[38][1] ),
    .B(_06489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06491_));
 sky130_fd_sc_hd__clkbuf_1 _13003_ (.A(_06491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01242_));
 sky130_fd_sc_hd__and2_1 _13004_ (.A(\sha256cu.m_pad_pars.block_512[38][2] ),
    .B(_06489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06492_));
 sky130_fd_sc_hd__clkbuf_1 _13005_ (.A(_06492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01243_));
 sky130_fd_sc_hd__and2_1 _13006_ (.A(\sha256cu.m_pad_pars.block_512[38][3] ),
    .B(_06489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06493_));
 sky130_fd_sc_hd__clkbuf_1 _13007_ (.A(_06493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01244_));
 sky130_fd_sc_hd__and2_1 _13008_ (.A(\sha256cu.m_pad_pars.block_512[38][4] ),
    .B(_06489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06494_));
 sky130_fd_sc_hd__clkbuf_1 _13009_ (.A(_06494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01245_));
 sky130_fd_sc_hd__and2_1 _13010_ (.A(\sha256cu.m_pad_pars.block_512[38][5] ),
    .B(_06489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06495_));
 sky130_fd_sc_hd__clkbuf_1 _13011_ (.A(_06495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01246_));
 sky130_fd_sc_hd__and2_1 _13012_ (.A(\sha256cu.m_pad_pars.block_512[38][6] ),
    .B(_06489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06496_));
 sky130_fd_sc_hd__clkbuf_1 _13013_ (.A(_06496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _13014_ (.A0(\sha256cu.m_pad_pars.block_512[38][7] ),
    .A1(_05085_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06497_));
 sky130_fd_sc_hd__clkbuf_1 _13015_ (.A(_06497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01248_));
 sky130_fd_sc_hd__o21ai_4 _13016_ (.A1(_04795_),
    .A2(_04970_),
    .B1(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06498_));
 sky130_fd_sc_hd__and2_1 _13017_ (.A(\sha256cu.m_pad_pars.block_512[39][0] ),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06499_));
 sky130_fd_sc_hd__clkbuf_1 _13018_ (.A(_06499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01249_));
 sky130_fd_sc_hd__and2_1 _13019_ (.A(\sha256cu.m_pad_pars.block_512[39][1] ),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06500_));
 sky130_fd_sc_hd__clkbuf_1 _13020_ (.A(_06500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01250_));
 sky130_fd_sc_hd__and2_1 _13021_ (.A(\sha256cu.m_pad_pars.block_512[39][2] ),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06501_));
 sky130_fd_sc_hd__clkbuf_1 _13022_ (.A(_06501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01251_));
 sky130_fd_sc_hd__and2_1 _13023_ (.A(\sha256cu.m_pad_pars.block_512[39][3] ),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06502_));
 sky130_fd_sc_hd__clkbuf_1 _13024_ (.A(_06502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01252_));
 sky130_fd_sc_hd__and2_1 _13025_ (.A(\sha256cu.m_pad_pars.block_512[39][4] ),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06503_));
 sky130_fd_sc_hd__clkbuf_1 _13026_ (.A(_06503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01253_));
 sky130_fd_sc_hd__and2_1 _13027_ (.A(\sha256cu.m_pad_pars.block_512[39][5] ),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06504_));
 sky130_fd_sc_hd__clkbuf_1 _13028_ (.A(_06504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01254_));
 sky130_fd_sc_hd__and2_1 _13029_ (.A(\sha256cu.m_pad_pars.block_512[39][6] ),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06505_));
 sky130_fd_sc_hd__clkbuf_1 _13030_ (.A(_06505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(\sha256cu.m_pad_pars.block_512[39][7] ),
    .A1(_04936_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06506_));
 sky130_fd_sc_hd__clkbuf_1 _13032_ (.A(_06506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01256_));
 sky130_fd_sc_hd__nand2_2 _13033_ (.A(_06270_),
    .B(_05319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06507_));
 sky130_fd_sc_hd__and2_1 _13034_ (.A(\sha256cu.m_pad_pars.block_512[40][0] ),
    .B(_06507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06508_));
 sky130_fd_sc_hd__clkbuf_1 _13035_ (.A(_06508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01257_));
 sky130_fd_sc_hd__and2_1 _13036_ (.A(\sha256cu.m_pad_pars.block_512[40][1] ),
    .B(_06507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06509_));
 sky130_fd_sc_hd__clkbuf_1 _13037_ (.A(_06509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01258_));
 sky130_fd_sc_hd__and2_1 _13038_ (.A(\sha256cu.m_pad_pars.block_512[40][2] ),
    .B(_06507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06510_));
 sky130_fd_sc_hd__clkbuf_1 _13039_ (.A(_06510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01259_));
 sky130_fd_sc_hd__and2_1 _13040_ (.A(\sha256cu.m_pad_pars.block_512[40][3] ),
    .B(_06507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06511_));
 sky130_fd_sc_hd__clkbuf_1 _13041_ (.A(_06511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01260_));
 sky130_fd_sc_hd__and2_1 _13042_ (.A(\sha256cu.m_pad_pars.block_512[40][4] ),
    .B(_06507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06512_));
 sky130_fd_sc_hd__clkbuf_1 _13043_ (.A(_06512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01261_));
 sky130_fd_sc_hd__and2_1 _13044_ (.A(\sha256cu.m_pad_pars.block_512[40][5] ),
    .B(_06507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06513_));
 sky130_fd_sc_hd__clkbuf_1 _13045_ (.A(_06513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01262_));
 sky130_fd_sc_hd__and2_1 _13046_ (.A(\sha256cu.m_pad_pars.block_512[40][6] ),
    .B(_06507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06514_));
 sky130_fd_sc_hd__clkbuf_1 _13047_ (.A(_06514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _13048_ (.A0(\sha256cu.m_pad_pars.block_512[40][7] ),
    .A1(_05400_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06515_));
 sky130_fd_sc_hd__clkbuf_1 _13049_ (.A(_06515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01264_));
 sky130_fd_sc_hd__or2_2 _13050_ (.A(_01986_),
    .B(_05131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06516_));
 sky130_fd_sc_hd__and2_1 _13051_ (.A(\sha256cu.m_pad_pars.block_512[41][0] ),
    .B(_06516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06517_));
 sky130_fd_sc_hd__clkbuf_1 _13052_ (.A(_06517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01265_));
 sky130_fd_sc_hd__and2_1 _13053_ (.A(\sha256cu.m_pad_pars.block_512[41][1] ),
    .B(_06516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06518_));
 sky130_fd_sc_hd__clkbuf_1 _13054_ (.A(_06518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01266_));
 sky130_fd_sc_hd__and2_1 _13055_ (.A(\sha256cu.m_pad_pars.block_512[41][2] ),
    .B(_06516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06519_));
 sky130_fd_sc_hd__clkbuf_1 _13056_ (.A(_06519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01267_));
 sky130_fd_sc_hd__and2_1 _13057_ (.A(\sha256cu.m_pad_pars.block_512[41][3] ),
    .B(_06516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06520_));
 sky130_fd_sc_hd__clkbuf_1 _13058_ (.A(_06520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01268_));
 sky130_fd_sc_hd__and2_1 _13059_ (.A(\sha256cu.m_pad_pars.block_512[41][4] ),
    .B(_06516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06521_));
 sky130_fd_sc_hd__clkbuf_1 _13060_ (.A(_06521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01269_));
 sky130_fd_sc_hd__and2_1 _13061_ (.A(\sha256cu.m_pad_pars.block_512[41][5] ),
    .B(_06516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06522_));
 sky130_fd_sc_hd__clkbuf_1 _13062_ (.A(_06522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01270_));
 sky130_fd_sc_hd__and2_1 _13063_ (.A(\sha256cu.m_pad_pars.block_512[41][6] ),
    .B(_06516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06523_));
 sky130_fd_sc_hd__clkbuf_1 _13064_ (.A(_06523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _13065_ (.A0(\sha256cu.m_pad_pars.block_512[41][7] ),
    .A1(_05232_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06524_));
 sky130_fd_sc_hd__clkbuf_1 _13066_ (.A(_06524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01272_));
 sky130_fd_sc_hd__or2_2 _13067_ (.A(_01986_),
    .B(_05000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06525_));
 sky130_fd_sc_hd__and2_1 _13068_ (.A(\sha256cu.m_pad_pars.block_512[42][0] ),
    .B(_06525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06526_));
 sky130_fd_sc_hd__clkbuf_1 _13069_ (.A(_06526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01273_));
 sky130_fd_sc_hd__and2_1 _13070_ (.A(\sha256cu.m_pad_pars.block_512[42][1] ),
    .B(_06525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06527_));
 sky130_fd_sc_hd__clkbuf_1 _13071_ (.A(_06527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01274_));
 sky130_fd_sc_hd__and2_1 _13072_ (.A(\sha256cu.m_pad_pars.block_512[42][2] ),
    .B(_06525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06528_));
 sky130_fd_sc_hd__clkbuf_1 _13073_ (.A(_06528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01275_));
 sky130_fd_sc_hd__and2_1 _13074_ (.A(\sha256cu.m_pad_pars.block_512[42][3] ),
    .B(_06525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06529_));
 sky130_fd_sc_hd__clkbuf_1 _13075_ (.A(_06529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01276_));
 sky130_fd_sc_hd__and2_1 _13076_ (.A(\sha256cu.m_pad_pars.block_512[42][4] ),
    .B(_06525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06530_));
 sky130_fd_sc_hd__clkbuf_1 _13077_ (.A(_06530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01277_));
 sky130_fd_sc_hd__and2_1 _13078_ (.A(\sha256cu.m_pad_pars.block_512[42][5] ),
    .B(_06525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06531_));
 sky130_fd_sc_hd__clkbuf_1 _13079_ (.A(_06531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01278_));
 sky130_fd_sc_hd__and2_1 _13080_ (.A(\sha256cu.m_pad_pars.block_512[42][6] ),
    .B(_06525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06532_));
 sky130_fd_sc_hd__clkbuf_1 _13081_ (.A(_06532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _13082_ (.A0(\sha256cu.m_pad_pars.block_512[42][7] ),
    .A1(_05087_),
    .S(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06533_));
 sky130_fd_sc_hd__clkbuf_1 _13083_ (.A(_06533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01280_));
 sky130_fd_sc_hd__or2_2 _13084_ (.A(_01986_),
    .B(_04803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06534_));
 sky130_fd_sc_hd__and2_1 _13085_ (.A(\sha256cu.m_pad_pars.block_512[43][0] ),
    .B(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06535_));
 sky130_fd_sc_hd__clkbuf_1 _13086_ (.A(_06535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01281_));
 sky130_fd_sc_hd__and2_1 _13087_ (.A(\sha256cu.m_pad_pars.block_512[43][1] ),
    .B(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06536_));
 sky130_fd_sc_hd__clkbuf_1 _13088_ (.A(_06536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01282_));
 sky130_fd_sc_hd__and2_1 _13089_ (.A(\sha256cu.m_pad_pars.block_512[43][2] ),
    .B(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06537_));
 sky130_fd_sc_hd__clkbuf_1 _13090_ (.A(_06537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01283_));
 sky130_fd_sc_hd__and2_1 _13091_ (.A(\sha256cu.m_pad_pars.block_512[43][3] ),
    .B(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06538_));
 sky130_fd_sc_hd__clkbuf_1 _13092_ (.A(_06538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01284_));
 sky130_fd_sc_hd__and2_1 _13093_ (.A(\sha256cu.m_pad_pars.block_512[43][4] ),
    .B(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06539_));
 sky130_fd_sc_hd__clkbuf_1 _13094_ (.A(_06539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01285_));
 sky130_fd_sc_hd__and2_1 _13095_ (.A(\sha256cu.m_pad_pars.block_512[43][5] ),
    .B(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06540_));
 sky130_fd_sc_hd__clkbuf_1 _13096_ (.A(_06540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01286_));
 sky130_fd_sc_hd__and2_1 _13097_ (.A(\sha256cu.m_pad_pars.block_512[43][6] ),
    .B(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06541_));
 sky130_fd_sc_hd__clkbuf_1 _13098_ (.A(_06541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01287_));
 sky130_fd_sc_hd__buf_4 _13099_ (.A(_01964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06542_));
 sky130_fd_sc_hd__mux2_1 _13100_ (.A0(\sha256cu.m_pad_pars.block_512[43][7] ),
    .A1(_04914_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06543_));
 sky130_fd_sc_hd__clkbuf_1 _13101_ (.A(_06543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01288_));
 sky130_fd_sc_hd__or3_2 _13102_ (.A(_02111_),
    .B(_04917_),
    .C(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06544_));
 sky130_fd_sc_hd__and2_1 _13103_ (.A(\sha256cu.m_pad_pars.block_512[44][0] ),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06545_));
 sky130_fd_sc_hd__clkbuf_1 _13104_ (.A(_06545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01289_));
 sky130_fd_sc_hd__and2_1 _13105_ (.A(\sha256cu.m_pad_pars.block_512[44][1] ),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06546_));
 sky130_fd_sc_hd__clkbuf_1 _13106_ (.A(_06546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01290_));
 sky130_fd_sc_hd__and2_1 _13107_ (.A(\sha256cu.m_pad_pars.block_512[44][2] ),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06547_));
 sky130_fd_sc_hd__clkbuf_1 _13108_ (.A(_06547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01291_));
 sky130_fd_sc_hd__and2_1 _13109_ (.A(\sha256cu.m_pad_pars.block_512[44][3] ),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06548_));
 sky130_fd_sc_hd__clkbuf_1 _13110_ (.A(_06548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01292_));
 sky130_fd_sc_hd__and2_1 _13111_ (.A(\sha256cu.m_pad_pars.block_512[44][4] ),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06549_));
 sky130_fd_sc_hd__clkbuf_1 _13112_ (.A(_06549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01293_));
 sky130_fd_sc_hd__and2_1 _13113_ (.A(\sha256cu.m_pad_pars.block_512[44][5] ),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06550_));
 sky130_fd_sc_hd__clkbuf_1 _13114_ (.A(_06550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01294_));
 sky130_fd_sc_hd__and2_1 _13115_ (.A(\sha256cu.m_pad_pars.block_512[44][6] ),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06551_));
 sky130_fd_sc_hd__clkbuf_1 _13116_ (.A(_06551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(\sha256cu.m_pad_pars.block_512[44][7] ),
    .A1(_05390_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06552_));
 sky130_fd_sc_hd__clkbuf_1 _13118_ (.A(_06552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01296_));
 sky130_fd_sc_hd__or3_2 _13119_ (.A(_02111_),
    .B(_04917_),
    .C(_05124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06553_));
 sky130_fd_sc_hd__and2_1 _13120_ (.A(\sha256cu.m_pad_pars.block_512[45][0] ),
    .B(_06553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06554_));
 sky130_fd_sc_hd__clkbuf_1 _13121_ (.A(_06554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01297_));
 sky130_fd_sc_hd__and2_1 _13122_ (.A(\sha256cu.m_pad_pars.block_512[45][1] ),
    .B(_06553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06555_));
 sky130_fd_sc_hd__clkbuf_1 _13123_ (.A(_06555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01298_));
 sky130_fd_sc_hd__and2_1 _13124_ (.A(\sha256cu.m_pad_pars.block_512[45][2] ),
    .B(_06553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06556_));
 sky130_fd_sc_hd__clkbuf_1 _13125_ (.A(_06556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01299_));
 sky130_fd_sc_hd__and2_1 _13126_ (.A(\sha256cu.m_pad_pars.block_512[45][3] ),
    .B(_06553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06557_));
 sky130_fd_sc_hd__clkbuf_1 _13127_ (.A(_06557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01300_));
 sky130_fd_sc_hd__and2_1 _13128_ (.A(\sha256cu.m_pad_pars.block_512[45][4] ),
    .B(_06553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06558_));
 sky130_fd_sc_hd__clkbuf_1 _13129_ (.A(_06558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01301_));
 sky130_fd_sc_hd__and2_1 _13130_ (.A(\sha256cu.m_pad_pars.block_512[45][5] ),
    .B(_06553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06559_));
 sky130_fd_sc_hd__clkbuf_1 _13131_ (.A(_06559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01302_));
 sky130_fd_sc_hd__and2_1 _13132_ (.A(\sha256cu.m_pad_pars.block_512[45][6] ),
    .B(_06553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06560_));
 sky130_fd_sc_hd__clkbuf_1 _13133_ (.A(_06560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(\sha256cu.m_pad_pars.block_512[45][7] ),
    .A1(_05256_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06561_));
 sky130_fd_sc_hd__clkbuf_1 _13135_ (.A(_06561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01304_));
 sky130_fd_sc_hd__or3_2 _13136_ (.A(_02111_),
    .B(_04917_),
    .C(_04975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06562_));
 sky130_fd_sc_hd__and2_1 _13137_ (.A(\sha256cu.m_pad_pars.block_512[46][0] ),
    .B(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06563_));
 sky130_fd_sc_hd__clkbuf_1 _13138_ (.A(_06563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01305_));
 sky130_fd_sc_hd__and2_1 _13139_ (.A(\sha256cu.m_pad_pars.block_512[46][1] ),
    .B(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06564_));
 sky130_fd_sc_hd__clkbuf_1 _13140_ (.A(_06564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01306_));
 sky130_fd_sc_hd__and2_1 _13141_ (.A(\sha256cu.m_pad_pars.block_512[46][2] ),
    .B(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06565_));
 sky130_fd_sc_hd__clkbuf_1 _13142_ (.A(_06565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01307_));
 sky130_fd_sc_hd__and2_1 _13143_ (.A(\sha256cu.m_pad_pars.block_512[46][3] ),
    .B(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06566_));
 sky130_fd_sc_hd__clkbuf_1 _13144_ (.A(_06566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01308_));
 sky130_fd_sc_hd__and2_1 _13145_ (.A(\sha256cu.m_pad_pars.block_512[46][4] ),
    .B(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06567_));
 sky130_fd_sc_hd__clkbuf_1 _13146_ (.A(_06567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01309_));
 sky130_fd_sc_hd__and2_1 _13147_ (.A(\sha256cu.m_pad_pars.block_512[46][5] ),
    .B(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06568_));
 sky130_fd_sc_hd__clkbuf_1 _13148_ (.A(_06568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01310_));
 sky130_fd_sc_hd__and2_1 _13149_ (.A(\sha256cu.m_pad_pars.block_512[46][6] ),
    .B(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06569_));
 sky130_fd_sc_hd__clkbuf_1 _13150_ (.A(_06569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(\sha256cu.m_pad_pars.block_512[46][7] ),
    .A1(_05113_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06570_));
 sky130_fd_sc_hd__clkbuf_1 _13152_ (.A(_06570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01312_));
 sky130_fd_sc_hd__or3_4 _13153_ (.A(_02111_),
    .B(_04705_),
    .C(_04820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06571_));
 sky130_fd_sc_hd__and2_1 _13154_ (.A(\sha256cu.m_pad_pars.block_512[47][0] ),
    .B(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06572_));
 sky130_fd_sc_hd__clkbuf_1 _13155_ (.A(_06572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01313_));
 sky130_fd_sc_hd__and2_1 _13156_ (.A(\sha256cu.m_pad_pars.block_512[47][1] ),
    .B(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06573_));
 sky130_fd_sc_hd__clkbuf_1 _13157_ (.A(_06573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01314_));
 sky130_fd_sc_hd__and2_1 _13158_ (.A(\sha256cu.m_pad_pars.block_512[47][2] ),
    .B(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06574_));
 sky130_fd_sc_hd__clkbuf_1 _13159_ (.A(_06574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01315_));
 sky130_fd_sc_hd__and2_1 _13160_ (.A(\sha256cu.m_pad_pars.block_512[47][3] ),
    .B(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06575_));
 sky130_fd_sc_hd__clkbuf_1 _13161_ (.A(_06575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01316_));
 sky130_fd_sc_hd__and2_1 _13162_ (.A(\sha256cu.m_pad_pars.block_512[47][4] ),
    .B(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06576_));
 sky130_fd_sc_hd__clkbuf_1 _13163_ (.A(_06576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01317_));
 sky130_fd_sc_hd__and2_1 _13164_ (.A(\sha256cu.m_pad_pars.block_512[47][5] ),
    .B(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06577_));
 sky130_fd_sc_hd__clkbuf_1 _13165_ (.A(_06577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01318_));
 sky130_fd_sc_hd__and2_1 _13166_ (.A(\sha256cu.m_pad_pars.block_512[47][6] ),
    .B(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06578_));
 sky130_fd_sc_hd__clkbuf_1 _13167_ (.A(_06578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _13168_ (.A0(\sha256cu.m_pad_pars.block_512[47][7] ),
    .A1(_04919_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06579_));
 sky130_fd_sc_hd__clkbuf_1 _13169_ (.A(_06579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01320_));
 sky130_fd_sc_hd__or3_2 _13170_ (.A(_02111_),
    .B(_04705_),
    .C(_05286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06580_));
 sky130_fd_sc_hd__and2_1 _13171_ (.A(\sha256cu.m_pad_pars.block_512[48][0] ),
    .B(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06581_));
 sky130_fd_sc_hd__clkbuf_1 _13172_ (.A(_06581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01321_));
 sky130_fd_sc_hd__and2_1 _13173_ (.A(\sha256cu.m_pad_pars.block_512[48][1] ),
    .B(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06582_));
 sky130_fd_sc_hd__clkbuf_1 _13174_ (.A(_06582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01322_));
 sky130_fd_sc_hd__and2_1 _13175_ (.A(\sha256cu.m_pad_pars.block_512[48][2] ),
    .B(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06583_));
 sky130_fd_sc_hd__clkbuf_1 _13176_ (.A(_06583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01323_));
 sky130_fd_sc_hd__and2_1 _13177_ (.A(\sha256cu.m_pad_pars.block_512[48][3] ),
    .B(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06584_));
 sky130_fd_sc_hd__clkbuf_1 _13178_ (.A(_06584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01324_));
 sky130_fd_sc_hd__and2_1 _13179_ (.A(\sha256cu.m_pad_pars.block_512[48][4] ),
    .B(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06585_));
 sky130_fd_sc_hd__clkbuf_1 _13180_ (.A(_06585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01325_));
 sky130_fd_sc_hd__and2_1 _13181_ (.A(\sha256cu.m_pad_pars.block_512[48][5] ),
    .B(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06586_));
 sky130_fd_sc_hd__clkbuf_1 _13182_ (.A(_06586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01326_));
 sky130_fd_sc_hd__and2_1 _13183_ (.A(\sha256cu.m_pad_pars.block_512[48][6] ),
    .B(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06587_));
 sky130_fd_sc_hd__clkbuf_1 _13184_ (.A(_06587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(\sha256cu.m_pad_pars.block_512[48][7] ),
    .A1(_05421_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06588_));
 sky130_fd_sc_hd__clkbuf_1 _13186_ (.A(_06588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01328_));
 sky130_fd_sc_hd__nor2_1 _13187_ (.A(_01952_),
    .B(_05136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06589_));
 sky130_fd_sc_hd__o21ai_4 _13188_ (.A1(_05269_),
    .A2(_06589_),
    .B1(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06590_));
 sky130_fd_sc_hd__and2_1 _13189_ (.A(\sha256cu.m_pad_pars.block_512[49][0] ),
    .B(_06590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06591_));
 sky130_fd_sc_hd__clkbuf_1 _13190_ (.A(_06591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01329_));
 sky130_fd_sc_hd__and2_1 _13191_ (.A(\sha256cu.m_pad_pars.block_512[49][1] ),
    .B(_06590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06592_));
 sky130_fd_sc_hd__clkbuf_1 _13192_ (.A(_06592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01330_));
 sky130_fd_sc_hd__and2_1 _13193_ (.A(\sha256cu.m_pad_pars.block_512[49][2] ),
    .B(_06590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06593_));
 sky130_fd_sc_hd__clkbuf_1 _13194_ (.A(_06593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01331_));
 sky130_fd_sc_hd__and2_1 _13195_ (.A(\sha256cu.m_pad_pars.block_512[49][3] ),
    .B(_06590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06594_));
 sky130_fd_sc_hd__clkbuf_1 _13196_ (.A(_06594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01332_));
 sky130_fd_sc_hd__and2_1 _13197_ (.A(\sha256cu.m_pad_pars.block_512[49][4] ),
    .B(_06590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06595_));
 sky130_fd_sc_hd__clkbuf_1 _13198_ (.A(_06595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01333_));
 sky130_fd_sc_hd__and2_1 _13199_ (.A(\sha256cu.m_pad_pars.block_512[49][5] ),
    .B(_06590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06596_));
 sky130_fd_sc_hd__clkbuf_1 _13200_ (.A(_06596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01334_));
 sky130_fd_sc_hd__and2_1 _13201_ (.A(\sha256cu.m_pad_pars.block_512[49][6] ),
    .B(_06590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06597_));
 sky130_fd_sc_hd__clkbuf_1 _13202_ (.A(_06597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _13203_ (.A0(\sha256cu.m_pad_pars.block_512[49][7] ),
    .A1(_05270_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06598_));
 sky130_fd_sc_hd__clkbuf_1 _13204_ (.A(_06598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01336_));
 sky130_fd_sc_hd__nand2_2 _13205_ (.A(_06270_),
    .B(_05006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06599_));
 sky130_fd_sc_hd__and2_1 _13206_ (.A(\sha256cu.m_pad_pars.block_512[50][0] ),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06600_));
 sky130_fd_sc_hd__clkbuf_1 _13207_ (.A(_06600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01337_));
 sky130_fd_sc_hd__and2_1 _13208_ (.A(\sha256cu.m_pad_pars.block_512[50][1] ),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06601_));
 sky130_fd_sc_hd__clkbuf_1 _13209_ (.A(_06601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01338_));
 sky130_fd_sc_hd__and2_1 _13210_ (.A(\sha256cu.m_pad_pars.block_512[50][2] ),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06602_));
 sky130_fd_sc_hd__clkbuf_1 _13211_ (.A(_06602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01339_));
 sky130_fd_sc_hd__and2_1 _13212_ (.A(\sha256cu.m_pad_pars.block_512[50][3] ),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06603_));
 sky130_fd_sc_hd__clkbuf_1 _13213_ (.A(_06603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01340_));
 sky130_fd_sc_hd__and2_1 _13214_ (.A(\sha256cu.m_pad_pars.block_512[50][4] ),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06604_));
 sky130_fd_sc_hd__clkbuf_1 _13215_ (.A(_06604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01341_));
 sky130_fd_sc_hd__and2_1 _13216_ (.A(\sha256cu.m_pad_pars.block_512[50][5] ),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06605_));
 sky130_fd_sc_hd__clkbuf_1 _13217_ (.A(_06605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01342_));
 sky130_fd_sc_hd__and2_1 _13218_ (.A(\sha256cu.m_pad_pars.block_512[50][6] ),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06606_));
 sky130_fd_sc_hd__clkbuf_1 _13219_ (.A(_06606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _13220_ (.A0(\sha256cu.m_pad_pars.block_512[50][7] ),
    .A1(_05109_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06607_));
 sky130_fd_sc_hd__clkbuf_1 _13221_ (.A(_06607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01344_));
 sky130_fd_sc_hd__o21ai_4 _13222_ (.A1(_04823_),
    .A2(_04825_),
    .B1(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06608_));
 sky130_fd_sc_hd__and2_1 _13223_ (.A(\sha256cu.m_pad_pars.block_512[51][0] ),
    .B(_06608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06609_));
 sky130_fd_sc_hd__clkbuf_1 _13224_ (.A(_06609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01345_));
 sky130_fd_sc_hd__and2_1 _13225_ (.A(\sha256cu.m_pad_pars.block_512[51][1] ),
    .B(_06608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06610_));
 sky130_fd_sc_hd__clkbuf_1 _13226_ (.A(_06610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01346_));
 sky130_fd_sc_hd__and2_1 _13227_ (.A(\sha256cu.m_pad_pars.block_512[51][2] ),
    .B(_06608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06611_));
 sky130_fd_sc_hd__clkbuf_1 _13228_ (.A(_06611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01347_));
 sky130_fd_sc_hd__and2_1 _13229_ (.A(\sha256cu.m_pad_pars.block_512[51][3] ),
    .B(_06608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06612_));
 sky130_fd_sc_hd__clkbuf_1 _13230_ (.A(_06612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01348_));
 sky130_fd_sc_hd__and2_1 _13231_ (.A(\sha256cu.m_pad_pars.block_512[51][4] ),
    .B(_06608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06613_));
 sky130_fd_sc_hd__clkbuf_1 _13232_ (.A(_06613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01349_));
 sky130_fd_sc_hd__and2_1 _13233_ (.A(\sha256cu.m_pad_pars.block_512[51][5] ),
    .B(_06608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06614_));
 sky130_fd_sc_hd__clkbuf_1 _13234_ (.A(_06614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01350_));
 sky130_fd_sc_hd__and2_1 _13235_ (.A(\sha256cu.m_pad_pars.block_512[51][6] ),
    .B(_06608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06615_));
 sky130_fd_sc_hd__clkbuf_1 _13236_ (.A(_06615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _13237_ (.A0(\sha256cu.m_pad_pars.block_512[51][7] ),
    .A1(_04932_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06616_));
 sky130_fd_sc_hd__clkbuf_1 _13238_ (.A(_06616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01352_));
 sky130_fd_sc_hd__nand2_2 _13239_ (.A(_06270_),
    .B(_05308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06617_));
 sky130_fd_sc_hd__and2_1 _13240_ (.A(\sha256cu.m_pad_pars.block_512[52][0] ),
    .B(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06618_));
 sky130_fd_sc_hd__clkbuf_1 _13241_ (.A(_06618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01353_));
 sky130_fd_sc_hd__and2_1 _13242_ (.A(\sha256cu.m_pad_pars.block_512[52][1] ),
    .B(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06619_));
 sky130_fd_sc_hd__clkbuf_1 _13243_ (.A(_06619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01354_));
 sky130_fd_sc_hd__and2_1 _13244_ (.A(\sha256cu.m_pad_pars.block_512[52][2] ),
    .B(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06620_));
 sky130_fd_sc_hd__clkbuf_1 _13245_ (.A(_06620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01355_));
 sky130_fd_sc_hd__and2_1 _13246_ (.A(\sha256cu.m_pad_pars.block_512[52][3] ),
    .B(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06621_));
 sky130_fd_sc_hd__clkbuf_1 _13247_ (.A(_06621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01356_));
 sky130_fd_sc_hd__and2_1 _13248_ (.A(\sha256cu.m_pad_pars.block_512[52][4] ),
    .B(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06622_));
 sky130_fd_sc_hd__clkbuf_1 _13249_ (.A(_06622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01357_));
 sky130_fd_sc_hd__and2_1 _13250_ (.A(\sha256cu.m_pad_pars.block_512[52][5] ),
    .B(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06623_));
 sky130_fd_sc_hd__clkbuf_1 _13251_ (.A(_06623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01358_));
 sky130_fd_sc_hd__and2_1 _13252_ (.A(\sha256cu.m_pad_pars.block_512[52][6] ),
    .B(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06624_));
 sky130_fd_sc_hd__clkbuf_1 _13253_ (.A(_06624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _13254_ (.A0(\sha256cu.m_pad_pars.block_512[52][7] ),
    .A1(_05415_),
    .S(_06542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06625_));
 sky130_fd_sc_hd__clkbuf_1 _13255_ (.A(_06625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01360_));
 sky130_fd_sc_hd__or4_4 _13256_ (.A(_02111_),
    .B(_01950_),
    .C(_04705_),
    .D(_05159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06626_));
 sky130_fd_sc_hd__and2_1 _13257_ (.A(\sha256cu.m_pad_pars.block_512[53][0] ),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06627_));
 sky130_fd_sc_hd__clkbuf_1 _13258_ (.A(_06627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01361_));
 sky130_fd_sc_hd__and2_1 _13259_ (.A(\sha256cu.m_pad_pars.block_512[53][1] ),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06628_));
 sky130_fd_sc_hd__clkbuf_1 _13260_ (.A(_06628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01362_));
 sky130_fd_sc_hd__and2_1 _13261_ (.A(\sha256cu.m_pad_pars.block_512[53][2] ),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06629_));
 sky130_fd_sc_hd__clkbuf_1 _13262_ (.A(_06629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01363_));
 sky130_fd_sc_hd__and2_1 _13263_ (.A(\sha256cu.m_pad_pars.block_512[53][3] ),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06630_));
 sky130_fd_sc_hd__clkbuf_1 _13264_ (.A(_06630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01364_));
 sky130_fd_sc_hd__and2_1 _13265_ (.A(\sha256cu.m_pad_pars.block_512[53][4] ),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06631_));
 sky130_fd_sc_hd__clkbuf_1 _13266_ (.A(_06631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01365_));
 sky130_fd_sc_hd__and2_1 _13267_ (.A(\sha256cu.m_pad_pars.block_512[53][5] ),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06632_));
 sky130_fd_sc_hd__clkbuf_1 _13268_ (.A(_06632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01366_));
 sky130_fd_sc_hd__and2_1 _13269_ (.A(\sha256cu.m_pad_pars.block_512[53][6] ),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06633_));
 sky130_fd_sc_hd__clkbuf_1 _13270_ (.A(_06633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _13271_ (.A0(\sha256cu.m_pad_pars.block_512[53][7] ),
    .A1(_05235_),
    .S(_01965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06634_));
 sky130_fd_sc_hd__clkbuf_1 _13272_ (.A(_06634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01368_));
 sky130_fd_sc_hd__a21o_2 _13273_ (.A1(_04979_),
    .A2(_04980_),
    .B1(_01912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06635_));
 sky130_fd_sc_hd__and2_1 _13274_ (.A(\sha256cu.m_pad_pars.block_512[54][0] ),
    .B(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06636_));
 sky130_fd_sc_hd__clkbuf_1 _13275_ (.A(_06636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01369_));
 sky130_fd_sc_hd__and2_1 _13276_ (.A(\sha256cu.m_pad_pars.block_512[54][1] ),
    .B(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06637_));
 sky130_fd_sc_hd__clkbuf_1 _13277_ (.A(_06637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01370_));
 sky130_fd_sc_hd__and2_1 _13278_ (.A(\sha256cu.m_pad_pars.block_512[54][2] ),
    .B(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06638_));
 sky130_fd_sc_hd__clkbuf_1 _13279_ (.A(_06638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01371_));
 sky130_fd_sc_hd__and2_1 _13280_ (.A(\sha256cu.m_pad_pars.block_512[54][3] ),
    .B(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06639_));
 sky130_fd_sc_hd__clkbuf_1 _13281_ (.A(_06639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01372_));
 sky130_fd_sc_hd__and2_1 _13282_ (.A(\sha256cu.m_pad_pars.block_512[54][4] ),
    .B(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06640_));
 sky130_fd_sc_hd__clkbuf_1 _13283_ (.A(_06640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01373_));
 sky130_fd_sc_hd__and2_1 _13284_ (.A(\sha256cu.m_pad_pars.block_512[54][5] ),
    .B(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06641_));
 sky130_fd_sc_hd__clkbuf_1 _13285_ (.A(_06641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01374_));
 sky130_fd_sc_hd__and2_1 _13286_ (.A(\sha256cu.m_pad_pars.block_512[54][6] ),
    .B(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06642_));
 sky130_fd_sc_hd__clkbuf_1 _13287_ (.A(_06642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _13288_ (.A0(\sha256cu.m_pad_pars.block_512[54][7] ),
    .A1(_05104_),
    .S(_01965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06643_));
 sky130_fd_sc_hd__clkbuf_1 _13289_ (.A(_06643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01376_));
 sky130_fd_sc_hd__or2_2 _13290_ (.A(_01986_),
    .B(_04832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06644_));
 sky130_fd_sc_hd__and2_1 _13291_ (.A(\sha256cu.m_pad_pars.block_512[55][0] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06645_));
 sky130_fd_sc_hd__clkbuf_1 _13292_ (.A(_06645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01377_));
 sky130_fd_sc_hd__and2_1 _13293_ (.A(\sha256cu.m_pad_pars.block_512[55][1] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06646_));
 sky130_fd_sc_hd__clkbuf_1 _13294_ (.A(_06646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01378_));
 sky130_fd_sc_hd__and2_1 _13295_ (.A(\sha256cu.m_pad_pars.block_512[55][2] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06647_));
 sky130_fd_sc_hd__clkbuf_1 _13296_ (.A(_06647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01379_));
 sky130_fd_sc_hd__and2_1 _13297_ (.A(\sha256cu.m_pad_pars.block_512[55][3] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06648_));
 sky130_fd_sc_hd__clkbuf_1 _13298_ (.A(_06648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01380_));
 sky130_fd_sc_hd__and2_1 _13299_ (.A(\sha256cu.m_pad_pars.block_512[55][4] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06649_));
 sky130_fd_sc_hd__clkbuf_1 _13300_ (.A(_06649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01381_));
 sky130_fd_sc_hd__and2_1 _13301_ (.A(\sha256cu.m_pad_pars.block_512[55][5] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06650_));
 sky130_fd_sc_hd__clkbuf_1 _13302_ (.A(_06650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01382_));
 sky130_fd_sc_hd__and2_1 _13303_ (.A(\sha256cu.m_pad_pars.block_512[55][6] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06651_));
 sky130_fd_sc_hd__clkbuf_1 _13304_ (.A(_06651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01383_));
 sky130_fd_sc_hd__and2_1 _13305_ (.A(\sha256cu.m_pad_pars.block_512[55][7] ),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06652_));
 sky130_fd_sc_hd__clkbuf_1 _13306_ (.A(_06652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01384_));
 sky130_fd_sc_hd__and2_1 _13307_ (.A(\sha256cu.m_pad_pars.block_512[56][0] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06653_));
 sky130_fd_sc_hd__clkbuf_1 _13308_ (.A(_06653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01385_));
 sky130_fd_sc_hd__and2_1 _13309_ (.A(\sha256cu.m_pad_pars.block_512[56][1] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06654_));
 sky130_fd_sc_hd__clkbuf_1 _13310_ (.A(_06654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01386_));
 sky130_fd_sc_hd__and2_1 _13311_ (.A(\sha256cu.m_pad_pars.block_512[56][2] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06655_));
 sky130_fd_sc_hd__clkbuf_1 _13312_ (.A(_06655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01387_));
 sky130_fd_sc_hd__and2_1 _13313_ (.A(\sha256cu.m_pad_pars.block_512[56][3] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06656_));
 sky130_fd_sc_hd__clkbuf_1 _13314_ (.A(_06656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01388_));
 sky130_fd_sc_hd__and2_1 _13315_ (.A(\sha256cu.m_pad_pars.block_512[56][4] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06657_));
 sky130_fd_sc_hd__clkbuf_1 _13316_ (.A(_06657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01389_));
 sky130_fd_sc_hd__and2_1 _13317_ (.A(\sha256cu.m_pad_pars.block_512[56][5] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06658_));
 sky130_fd_sc_hd__clkbuf_1 _13318_ (.A(_06658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01390_));
 sky130_fd_sc_hd__and2_1 _13319_ (.A(\sha256cu.m_pad_pars.block_512[56][6] ),
    .B(_01924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06659_));
 sky130_fd_sc_hd__clkbuf_1 _13320_ (.A(_06659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01391_));
 sky130_fd_sc_hd__buf_2 _13321_ (.A(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06660_));
 sky130_fd_sc_hd__and2_1 _13322_ (.A(\sha256cu.m_pad_pars.block_512[56][7] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06661_));
 sky130_fd_sc_hd__clkbuf_1 _13323_ (.A(_06661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01392_));
 sky130_fd_sc_hd__and2_1 _13324_ (.A(\sha256cu.m_pad_pars.block_512[57][0] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06662_));
 sky130_fd_sc_hd__clkbuf_1 _13325_ (.A(_06662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01393_));
 sky130_fd_sc_hd__and2_1 _13326_ (.A(\sha256cu.m_pad_pars.block_512[57][1] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06663_));
 sky130_fd_sc_hd__clkbuf_1 _13327_ (.A(_06663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01394_));
 sky130_fd_sc_hd__and2_1 _13328_ (.A(\sha256cu.m_pad_pars.block_512[57][2] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06664_));
 sky130_fd_sc_hd__clkbuf_1 _13329_ (.A(_06664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01395_));
 sky130_fd_sc_hd__and2_1 _13330_ (.A(\sha256cu.m_pad_pars.block_512[57][3] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06665_));
 sky130_fd_sc_hd__clkbuf_1 _13331_ (.A(_06665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01396_));
 sky130_fd_sc_hd__and2_1 _13332_ (.A(\sha256cu.m_pad_pars.block_512[57][4] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06666_));
 sky130_fd_sc_hd__clkbuf_1 _13333_ (.A(_06666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01397_));
 sky130_fd_sc_hd__and2_1 _13334_ (.A(\sha256cu.m_pad_pars.block_512[57][5] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06667_));
 sky130_fd_sc_hd__clkbuf_1 _13335_ (.A(_06667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01398_));
 sky130_fd_sc_hd__and2_1 _13336_ (.A(\sha256cu.m_pad_pars.block_512[57][6] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06668_));
 sky130_fd_sc_hd__clkbuf_1 _13337_ (.A(_06668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01399_));
 sky130_fd_sc_hd__and2_1 _13338_ (.A(\sha256cu.m_pad_pars.block_512[57][7] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06669_));
 sky130_fd_sc_hd__clkbuf_1 _13339_ (.A(_06669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01400_));
 sky130_fd_sc_hd__and2_1 _13340_ (.A(\sha256cu.m_pad_pars.block_512[58][0] ),
    .B(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06670_));
 sky130_fd_sc_hd__clkbuf_1 _13341_ (.A(_06670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01401_));
 sky130_fd_sc_hd__clkbuf_4 _13342_ (.A(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06671_));
 sky130_fd_sc_hd__and2_1 _13343_ (.A(\sha256cu.m_pad_pars.block_512[58][1] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06672_));
 sky130_fd_sc_hd__clkbuf_1 _13344_ (.A(_06672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01402_));
 sky130_fd_sc_hd__and2_1 _13345_ (.A(\sha256cu.m_pad_pars.block_512[58][2] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06673_));
 sky130_fd_sc_hd__clkbuf_1 _13346_ (.A(_06673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01403_));
 sky130_fd_sc_hd__and2_1 _13347_ (.A(\sha256cu.m_pad_pars.block_512[58][3] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06674_));
 sky130_fd_sc_hd__clkbuf_1 _13348_ (.A(_06674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01404_));
 sky130_fd_sc_hd__and2_1 _13349_ (.A(\sha256cu.m_pad_pars.block_512[58][4] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06675_));
 sky130_fd_sc_hd__clkbuf_1 _13350_ (.A(_06675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01405_));
 sky130_fd_sc_hd__and2_1 _13351_ (.A(\sha256cu.m_pad_pars.block_512[58][5] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06676_));
 sky130_fd_sc_hd__clkbuf_1 _13352_ (.A(_06676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01406_));
 sky130_fd_sc_hd__and2_1 _13353_ (.A(\sha256cu.m_pad_pars.block_512[58][6] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06677_));
 sky130_fd_sc_hd__clkbuf_1 _13354_ (.A(_06677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01407_));
 sky130_fd_sc_hd__and2_1 _13355_ (.A(\sha256cu.m_pad_pars.block_512[58][7] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06678_));
 sky130_fd_sc_hd__clkbuf_1 _13356_ (.A(_06678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01408_));
 sky130_fd_sc_hd__and2_1 _13357_ (.A(\sha256cu.m_pad_pars.block_512[59][0] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06679_));
 sky130_fd_sc_hd__clkbuf_1 _13358_ (.A(_06679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01409_));
 sky130_fd_sc_hd__and2_1 _13359_ (.A(\sha256cu.m_pad_pars.block_512[59][1] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06680_));
 sky130_fd_sc_hd__clkbuf_1 _13360_ (.A(_06680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01410_));
 sky130_fd_sc_hd__and2_1 _13361_ (.A(\sha256cu.m_pad_pars.block_512[59][2] ),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06681_));
 sky130_fd_sc_hd__clkbuf_1 _13362_ (.A(_06681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01411_));
 sky130_fd_sc_hd__buf_2 _13363_ (.A(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06682_));
 sky130_fd_sc_hd__and2_1 _13364_ (.A(\sha256cu.m_pad_pars.block_512[59][3] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06683_));
 sky130_fd_sc_hd__clkbuf_1 _13365_ (.A(_06683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01412_));
 sky130_fd_sc_hd__and2_1 _13366_ (.A(\sha256cu.m_pad_pars.block_512[59][4] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06684_));
 sky130_fd_sc_hd__clkbuf_1 _13367_ (.A(_06684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01413_));
 sky130_fd_sc_hd__and2_1 _13368_ (.A(\sha256cu.m_pad_pars.block_512[59][5] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06685_));
 sky130_fd_sc_hd__clkbuf_1 _13369_ (.A(_06685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01414_));
 sky130_fd_sc_hd__and2_1 _13370_ (.A(\sha256cu.m_pad_pars.block_512[59][6] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06686_));
 sky130_fd_sc_hd__clkbuf_1 _13371_ (.A(_06686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01415_));
 sky130_fd_sc_hd__and2_1 _13372_ (.A(\sha256cu.m_pad_pars.block_512[59][7] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06687_));
 sky130_fd_sc_hd__clkbuf_1 _13373_ (.A(_06687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01416_));
 sky130_fd_sc_hd__and2_1 _13374_ (.A(\sha256cu.m_pad_pars.block_512[60][0] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06688_));
 sky130_fd_sc_hd__clkbuf_1 _13375_ (.A(_06688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01417_));
 sky130_fd_sc_hd__and2_1 _13376_ (.A(\sha256cu.m_pad_pars.block_512[60][1] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06689_));
 sky130_fd_sc_hd__clkbuf_1 _13377_ (.A(_06689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01418_));
 sky130_fd_sc_hd__and2_1 _13378_ (.A(\sha256cu.m_pad_pars.block_512[60][2] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06690_));
 sky130_fd_sc_hd__clkbuf_1 _13379_ (.A(_06690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01419_));
 sky130_fd_sc_hd__and2_1 _13380_ (.A(\sha256cu.m_pad_pars.block_512[60][3] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06691_));
 sky130_fd_sc_hd__clkbuf_1 _13381_ (.A(_06691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01420_));
 sky130_fd_sc_hd__and2_1 _13382_ (.A(\sha256cu.m_pad_pars.block_512[60][4] ),
    .B(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06692_));
 sky130_fd_sc_hd__clkbuf_1 _13383_ (.A(_06692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01421_));
 sky130_fd_sc_hd__buf_2 _13384_ (.A(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06693_));
 sky130_fd_sc_hd__and2_1 _13385_ (.A(\sha256cu.m_pad_pars.block_512[60][5] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06694_));
 sky130_fd_sc_hd__clkbuf_1 _13386_ (.A(_06694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01422_));
 sky130_fd_sc_hd__and2_1 _13387_ (.A(\sha256cu.m_pad_pars.block_512[60][6] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06695_));
 sky130_fd_sc_hd__clkbuf_1 _13388_ (.A(_06695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01423_));
 sky130_fd_sc_hd__and2_1 _13389_ (.A(\sha256cu.m_pad_pars.block_512[60][7] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06696_));
 sky130_fd_sc_hd__clkbuf_1 _13390_ (.A(_06696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01424_));
 sky130_fd_sc_hd__and2_1 _13391_ (.A(\sha256cu.m_pad_pars.block_512[61][0] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06697_));
 sky130_fd_sc_hd__clkbuf_1 _13392_ (.A(_06697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01425_));
 sky130_fd_sc_hd__and2_1 _13393_ (.A(\sha256cu.m_pad_pars.block_512[61][1] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06698_));
 sky130_fd_sc_hd__clkbuf_1 _13394_ (.A(_06698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01426_));
 sky130_fd_sc_hd__and2_1 _13395_ (.A(\sha256cu.m_pad_pars.block_512[61][2] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06699_));
 sky130_fd_sc_hd__clkbuf_1 _13396_ (.A(_06699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01427_));
 sky130_fd_sc_hd__and2_1 _13397_ (.A(\sha256cu.m_pad_pars.block_512[61][3] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06700_));
 sky130_fd_sc_hd__clkbuf_1 _13398_ (.A(_06700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01428_));
 sky130_fd_sc_hd__and2_1 _13399_ (.A(\sha256cu.m_pad_pars.block_512[61][4] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06701_));
 sky130_fd_sc_hd__clkbuf_1 _13400_ (.A(_06701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01429_));
 sky130_fd_sc_hd__and2_1 _13401_ (.A(\sha256cu.m_pad_pars.block_512[61][5] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_1 _13402_ (.A(_06702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01430_));
 sky130_fd_sc_hd__and2_1 _13403_ (.A(\sha256cu.m_pad_pars.block_512[61][6] ),
    .B(_06693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06703_));
 sky130_fd_sc_hd__clkbuf_1 _13404_ (.A(_06703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01431_));
 sky130_fd_sc_hd__and2_1 _13405_ (.A(\sha256cu.m_pad_pars.block_512[61][7] ),
    .B(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06704_));
 sky130_fd_sc_hd__clkbuf_1 _13406_ (.A(_06704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _13407_ (.A0(\sha256cu.m_pad_pars.m_size[8] ),
    .A1(\sha256cu.m_pad_pars.block_512[62][0] ),
    .S(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06705_));
 sky130_fd_sc_hd__clkbuf_1 _13408_ (.A(_06705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _13409_ (.A0(\sha256cu.m_pad_pars.m_size[9] ),
    .A1(\sha256cu.m_pad_pars.block_512[62][1] ),
    .S(_01923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06706_));
 sky130_fd_sc_hd__clkbuf_1 _13410_ (.A(_06706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01434_));
 sky130_fd_sc_hd__and2_1 _13411_ (.A(\sha256cu.m_pad_pars.block_512[62][2] ),
    .B(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06707_));
 sky130_fd_sc_hd__clkbuf_1 _13412_ (.A(_06707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01435_));
 sky130_fd_sc_hd__and2_1 _13413_ (.A(\sha256cu.m_pad_pars.block_512[62][3] ),
    .B(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06708_));
 sky130_fd_sc_hd__clkbuf_1 _13414_ (.A(_06708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01436_));
 sky130_fd_sc_hd__and2_1 _13415_ (.A(\sha256cu.m_pad_pars.block_512[62][4] ),
    .B(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06709_));
 sky130_fd_sc_hd__clkbuf_1 _13416_ (.A(_06709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01437_));
 sky130_fd_sc_hd__and2_1 _13417_ (.A(\sha256cu.m_pad_pars.block_512[62][5] ),
    .B(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06710_));
 sky130_fd_sc_hd__clkbuf_1 _13418_ (.A(_06710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01438_));
 sky130_fd_sc_hd__and2_1 _13419_ (.A(\sha256cu.m_pad_pars.block_512[62][6] ),
    .B(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06711_));
 sky130_fd_sc_hd__clkbuf_1 _13420_ (.A(_06711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01439_));
 sky130_fd_sc_hd__and2_1 _13421_ (.A(\sha256cu.m_pad_pars.block_512[62][7] ),
    .B(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06712_));
 sky130_fd_sc_hd__clkbuf_1 _13422_ (.A(_06712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01440_));
 sky130_fd_sc_hd__nor2_4 _13423_ (.A(\sha256cu.temp_case ),
    .B(_04177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06713_));
 sky130_fd_sc_hd__clkbuf_4 _13424_ (.A(_06713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06714_));
 sky130_fd_sc_hd__or2_1 _13425_ (.A(\sha256cu.temp_case ),
    .B(_04177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06715_));
 sky130_fd_sc_hd__clkbuf_2 _13426_ (.A(_06715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06716_));
 sky130_fd_sc_hd__nand2_2 _13427_ (.A(\sha256cu.iter_processing.padding_done ),
    .B(_06716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06717_));
 sky130_fd_sc_hd__nor2_4 _13428_ (.A(\sha256cu.counter_iteration[6] ),
    .B(_06717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06718_));
 sky130_fd_sc_hd__clkbuf_4 _13429_ (.A(_06718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06719_));
 sky130_fd_sc_hd__a22o_1 _13430_ (.A1(\sha256cu.K[0] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06720_));
 sky130_fd_sc_hd__and2_1 _13431_ (.A(_03288_),
    .B(_06720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06721_));
 sky130_fd_sc_hd__clkbuf_1 _13432_ (.A(_06721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01441_));
 sky130_fd_sc_hd__a22o_1 _13433_ (.A1(\sha256cu.K[1] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06722_));
 sky130_fd_sc_hd__and2_1 _13434_ (.A(_03288_),
    .B(_06722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06723_));
 sky130_fd_sc_hd__clkbuf_1 _13435_ (.A(_06723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01442_));
 sky130_fd_sc_hd__a22o_1 _13436_ (.A1(\sha256cu.K[2] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06724_));
 sky130_fd_sc_hd__and2_1 _13437_ (.A(_03288_),
    .B(_06724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06725_));
 sky130_fd_sc_hd__clkbuf_1 _13438_ (.A(_06725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01443_));
 sky130_fd_sc_hd__clkbuf_4 _13439_ (.A(_06716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06726_));
 sky130_fd_sc_hd__buf_2 _13440_ (.A(_06717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06727_));
 sky130_fd_sc_hd__and2b_1 _13441_ (.A_N(_04188_),
    .B(_00061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06728_));
 sky130_fd_sc_hd__o221a_1 _13442_ (.A1(\sha256cu.K[3] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06728_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01444_));
 sky130_fd_sc_hd__and2b_1 _13443_ (.A_N(_04188_),
    .B(_00062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06729_));
 sky130_fd_sc_hd__o221a_1 _13444_ (.A1(\sha256cu.K[4] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06729_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01445_));
 sky130_fd_sc_hd__buf_2 _13445_ (.A(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06730_));
 sky130_fd_sc_hd__a22o_1 _13446_ (.A1(\sha256cu.K[5] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06731_));
 sky130_fd_sc_hd__and2_1 _13447_ (.A(_06730_),
    .B(_06731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06732_));
 sky130_fd_sc_hd__clkbuf_1 _13448_ (.A(_06732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01446_));
 sky130_fd_sc_hd__a22o_1 _13449_ (.A1(\sha256cu.K[6] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06733_));
 sky130_fd_sc_hd__and2_1 _13450_ (.A(_06730_),
    .B(_06733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06734_));
 sky130_fd_sc_hd__clkbuf_1 _13451_ (.A(_06734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01447_));
 sky130_fd_sc_hd__and2b_1 _13452_ (.A_N(_04188_),
    .B(_00065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06735_));
 sky130_fd_sc_hd__o221a_1 _13453_ (.A1(\sha256cu.K[7] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06735_),
    .C1(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01448_));
 sky130_fd_sc_hd__and2b_1 _13454_ (.A_N(_04188_),
    .B(_00066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06736_));
 sky130_fd_sc_hd__buf_2 _13455_ (.A(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06737_));
 sky130_fd_sc_hd__o221a_1 _13456_ (.A1(\sha256cu.K[8] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06736_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01449_));
 sky130_fd_sc_hd__and2b_1 _13457_ (.A_N(_04188_),
    .B(_00067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06738_));
 sky130_fd_sc_hd__o221a_1 _13458_ (.A1(\sha256cu.K[9] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06738_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01450_));
 sky130_fd_sc_hd__and2b_1 _13459_ (.A_N(_04188_),
    .B(_00037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06739_));
 sky130_fd_sc_hd__o221a_1 _13460_ (.A1(\sha256cu.K[10] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06739_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01451_));
 sky130_fd_sc_hd__and2b_1 _13461_ (.A_N(_04188_),
    .B(_00038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06740_));
 sky130_fd_sc_hd__o221a_1 _13462_ (.A1(\sha256cu.K[11] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06740_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01452_));
 sky130_fd_sc_hd__a22o_1 _13463_ (.A1(\sha256cu.K[12] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06741_));
 sky130_fd_sc_hd__and2_1 _13464_ (.A(_06730_),
    .B(_06741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06742_));
 sky130_fd_sc_hd__clkbuf_1 _13465_ (.A(_06742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01453_));
 sky130_fd_sc_hd__and2b_1 _13466_ (.A_N(_04188_),
    .B(_00040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06743_));
 sky130_fd_sc_hd__o221a_1 _13467_ (.A1(\sha256cu.K[13] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06743_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01454_));
 sky130_fd_sc_hd__a22o_1 _13468_ (.A1(\sha256cu.K[14] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06744_));
 sky130_fd_sc_hd__and2_1 _13469_ (.A(_06730_),
    .B(_06744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06745_));
 sky130_fd_sc_hd__clkbuf_1 _13470_ (.A(_06745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01455_));
 sky130_fd_sc_hd__a22o_1 _13471_ (.A1(\sha256cu.K[15] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06746_));
 sky130_fd_sc_hd__and2_1 _13472_ (.A(_06730_),
    .B(_06746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06747_));
 sky130_fd_sc_hd__clkbuf_1 _13473_ (.A(_06747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01456_));
 sky130_fd_sc_hd__a22o_1 _13474_ (.A1(\sha256cu.K[16] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06748_));
 sky130_fd_sc_hd__and2_1 _13475_ (.A(_06730_),
    .B(_06748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06749_));
 sky130_fd_sc_hd__clkbuf_1 _13476_ (.A(_06749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01457_));
 sky130_fd_sc_hd__and2b_1 _13477_ (.A_N(_04188_),
    .B(_00044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06750_));
 sky130_fd_sc_hd__o221a_1 _13478_ (.A1(\sha256cu.K[17] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06750_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01458_));
 sky130_fd_sc_hd__a22o_1 _13479_ (.A1(\sha256cu.K[18] ),
    .A2(_06714_),
    .B1(_06719_),
    .B2(_00045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06751_));
 sky130_fd_sc_hd__and2_1 _13480_ (.A(_06730_),
    .B(_06751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06752_));
 sky130_fd_sc_hd__clkbuf_1 _13481_ (.A(_06752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01459_));
 sky130_fd_sc_hd__and2b_1 _13482_ (.A_N(\sha256cu.counter_iteration[6] ),
    .B(_00046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06753_));
 sky130_fd_sc_hd__o221a_1 _13483_ (.A1(\sha256cu.K[19] ),
    .A2(_06726_),
    .B1(_06727_),
    .B2(_06753_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01460_));
 sky130_fd_sc_hd__a22o_1 _13484_ (.A1(\sha256cu.K[20] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06754_));
 sky130_fd_sc_hd__and2_1 _13485_ (.A(_06730_),
    .B(_06754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06755_));
 sky130_fd_sc_hd__clkbuf_1 _13486_ (.A(_06755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01461_));
 sky130_fd_sc_hd__a22o_1 _13487_ (.A1(\sha256cu.K[21] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06756_));
 sky130_fd_sc_hd__and2_1 _13488_ (.A(_06730_),
    .B(_06756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06757_));
 sky130_fd_sc_hd__clkbuf_1 _13489_ (.A(_06757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01462_));
 sky130_fd_sc_hd__a22o_1 _13490_ (.A1(\sha256cu.K[22] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06758_));
 sky130_fd_sc_hd__and2_1 _13491_ (.A(_06730_),
    .B(_06758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06759_));
 sky130_fd_sc_hd__clkbuf_1 _13492_ (.A(_06759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01463_));
 sky130_fd_sc_hd__and2b_1 _13493_ (.A_N(\sha256cu.counter_iteration[6] ),
    .B(_00051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06760_));
 sky130_fd_sc_hd__o221a_1 _13494_ (.A1(\sha256cu.K[23] ),
    .A2(_06716_),
    .B1(_06717_),
    .B2(_06760_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01464_));
 sky130_fd_sc_hd__a22o_1 _13495_ (.A1(\sha256cu.K[24] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06761_));
 sky130_fd_sc_hd__and2_1 _13496_ (.A(_01975_),
    .B(_06761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06762_));
 sky130_fd_sc_hd__clkbuf_1 _13497_ (.A(_06762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01465_));
 sky130_fd_sc_hd__and2b_1 _13498_ (.A_N(\sha256cu.counter_iteration[6] ),
    .B(_00053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06763_));
 sky130_fd_sc_hd__o221a_1 _13499_ (.A1(\sha256cu.K[25] ),
    .A2(_06716_),
    .B1(_06717_),
    .B2(_06763_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01466_));
 sky130_fd_sc_hd__a22o_1 _13500_ (.A1(\sha256cu.K[26] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06764_));
 sky130_fd_sc_hd__and2_1 _13501_ (.A(_01975_),
    .B(_06764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06765_));
 sky130_fd_sc_hd__clkbuf_1 _13502_ (.A(_06765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01467_));
 sky130_fd_sc_hd__a22o_1 _13503_ (.A1(\sha256cu.K[27] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06766_));
 sky130_fd_sc_hd__and2_1 _13504_ (.A(_01975_),
    .B(_06766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06767_));
 sky130_fd_sc_hd__clkbuf_1 _13505_ (.A(_06767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01468_));
 sky130_fd_sc_hd__a22o_1 _13506_ (.A1(\sha256cu.K[28] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06768_));
 sky130_fd_sc_hd__and2_1 _13507_ (.A(_01975_),
    .B(_06768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06769_));
 sky130_fd_sc_hd__clkbuf_1 _13508_ (.A(_06769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01469_));
 sky130_fd_sc_hd__a22o_1 _13509_ (.A1(\sha256cu.K[29] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06770_));
 sky130_fd_sc_hd__and2_1 _13510_ (.A(_01975_),
    .B(_06770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06771_));
 sky130_fd_sc_hd__clkbuf_1 _13511_ (.A(_06771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01470_));
 sky130_fd_sc_hd__and2b_1 _13512_ (.A_N(\sha256cu.counter_iteration[6] ),
    .B(_00059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06772_));
 sky130_fd_sc_hd__o221a_1 _13513_ (.A1(\sha256cu.K[30] ),
    .A2(_06716_),
    .B1(_06717_),
    .B2(_06772_),
    .C1(_06737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01471_));
 sky130_fd_sc_hd__a22o_1 _13514_ (.A1(\sha256cu.K[31] ),
    .A2(_06713_),
    .B1(_06718_),
    .B2(_00060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06773_));
 sky130_fd_sc_hd__and2_1 _13515_ (.A(_01975_),
    .B(_06773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06774_));
 sky130_fd_sc_hd__clkbuf_1 _13516_ (.A(_06774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01472_));
 sky130_fd_sc_hd__o21a_1 _13517_ (.A1(\sha256cu.temp_case ),
    .A2(\sha256cu.iter_processing.padding_done ),
    .B1(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01473_));
 sky130_fd_sc_hd__dfxtp_1 _13518_ (.CLK(clknet_leaf_108_clk),
    .D(_00068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.byte_stop ));
 sky130_fd_sc_hd__dfxtp_2 _13519_ (.CLK(clknet_leaf_79_clk),
    .D(_00069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net258));
 sky130_fd_sc_hd__dfxtp_1 _13520_ (.CLK(clknet_leaf_109_clk),
    .D(_00070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net259));
 sky130_fd_sc_hd__dfxtp_4 _13521_ (.CLK(clknet_leaf_79_clk),
    .D(_00071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.rst ));
 sky130_fd_sc_hd__dfxtp_1 _13522_ (.CLK(clknet_leaf_124_clk),
    .D(_00072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13523_ (.CLK(clknet_leaf_125_clk),
    .D(_00073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13524_ (.CLK(clknet_leaf_1_clk),
    .D(_00074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13525_ (.CLK(clknet_leaf_2_clk),
    .D(_00075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13526_ (.CLK(clknet_leaf_124_clk),
    .D(_00076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13527_ (.CLK(clknet_leaf_124_clk),
    .D(_00077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13528_ (.CLK(clknet_leaf_2_clk),
    .D(_00078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13529_ (.CLK(clknet_leaf_123_clk),
    .D(_00079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[63][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13530_ (.CLK(clknet_leaf_108_clk),
    .D(_00080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.byte_rdy ));
 sky130_fd_sc_hd__dfxtp_2 _13531_ (.CLK(clknet_leaf_107_clk),
    .D(_00081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13532_ (.CLK(clknet_leaf_107_clk),
    .D(_00082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13533_ (.CLK(clknet_leaf_107_clk),
    .D(_00083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13534_ (.CLK(clknet_leaf_103_clk),
    .D(_00084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13535_ (.CLK(clknet_leaf_109_clk),
    .D(_00032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13536_ (.CLK(clknet_leaf_79_clk),
    .D(_00033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13537_ (.CLK(clknet_leaf_109_clk),
    .D(_00034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13538_ (.CLK(clknet_leaf_109_clk),
    .D(_00035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13539_ (.CLK(clknet_leaf_112_clk),
    .D(_00085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13540_ (.CLK(clknet_leaf_112_clk),
    .D(_00086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out0[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13541_ (.CLK(clknet_leaf_117_clk),
    .D(_00087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13542_ (.CLK(clknet_leaf_117_clk),
    .D(_00088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13543_ (.CLK(clknet_leaf_107_clk),
    .D(_00089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13544_ (.CLK(clknet_leaf_105_clk),
    .D(_00090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.temp_if ));
 sky130_fd_sc_hd__dfxtp_1 _13545_ (.CLK(clknet_leaf_79_clk),
    .D(_00091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(Hash_Digest));
 sky130_fd_sc_hd__dfxtp_1 _13546_ (.CLK(clknet_leaf_105_clk),
    .D(_00092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.temp_delay ));
 sky130_fd_sc_hd__dfxtp_1 _13547_ (.CLK(clknet_leaf_79_clk),
    .D(_00093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.H7[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13548_ (.CLK(clknet_leaf_80_clk),
    .D(_00094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.temp_case ));
 sky130_fd_sc_hd__dfxtp_2 _13549_ (.CLK(clknet_leaf_74_clk),
    .D(_00095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[0] ));
 sky130_fd_sc_hd__dfxtp_4 _13550_ (.CLK(clknet_leaf_75_clk),
    .D(_00096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[1] ));
 sky130_fd_sc_hd__dfxtp_4 _13551_ (.CLK(clknet_leaf_73_clk),
    .D(_00097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[2] ));
 sky130_fd_sc_hd__dfxtp_4 _13552_ (.CLK(clknet_leaf_51_clk),
    .D(_00098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[3] ));
 sky130_fd_sc_hd__dfxtp_4 _13553_ (.CLK(clknet_leaf_51_clk),
    .D(_00099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[4] ));
 sky130_fd_sc_hd__dfxtp_4 _13554_ (.CLK(clknet_leaf_51_clk),
    .D(_00100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[5] ));
 sky130_fd_sc_hd__dfxtp_4 _13555_ (.CLK(clknet_leaf_51_clk),
    .D(_00101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[6] ));
 sky130_fd_sc_hd__dfxtp_4 _13556_ (.CLK(clknet_leaf_59_clk),
    .D(_00102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[7] ));
 sky130_fd_sc_hd__dfxtp_4 _13557_ (.CLK(clknet_leaf_61_clk),
    .D(_00103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[8] ));
 sky130_fd_sc_hd__dfxtp_4 _13558_ (.CLK(clknet_leaf_65_clk),
    .D(_00104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[9] ));
 sky130_fd_sc_hd__dfxtp_4 _13559_ (.CLK(clknet_leaf_63_clk),
    .D(_00105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[10] ));
 sky130_fd_sc_hd__dfxtp_4 _13560_ (.CLK(clknet_leaf_68_clk),
    .D(_00106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13561_ (.CLK(clknet_leaf_64_clk),
    .D(_00107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13562_ (.CLK(clknet_leaf_64_clk),
    .D(_00108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[13] ));
 sky130_fd_sc_hd__dfxtp_4 _13563_ (.CLK(clknet_leaf_65_clk),
    .D(_00109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13564_ (.CLK(clknet_leaf_64_clk),
    .D(_00110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13565_ (.CLK(clknet_leaf_69_clk),
    .D(_00111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13566_ (.CLK(clknet_leaf_69_clk),
    .D(_00112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13567_ (.CLK(clknet_leaf_69_clk),
    .D(_00113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13568_ (.CLK(clknet_leaf_69_clk),
    .D(_00114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13569_ (.CLK(clknet_leaf_85_clk),
    .D(_00115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[20] ));
 sky130_fd_sc_hd__dfxtp_4 _13570_ (.CLK(clknet_leaf_85_clk),
    .D(_00116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13571_ (.CLK(clknet_leaf_86_clk),
    .D(_00117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[22] ));
 sky130_fd_sc_hd__dfxtp_4 _13572_ (.CLK(clknet_leaf_85_clk),
    .D(_00118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13573_ (.CLK(clknet_leaf_86_clk),
    .D(_00119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[24] ));
 sky130_fd_sc_hd__dfxtp_4 _13574_ (.CLK(clknet_leaf_85_clk),
    .D(_00120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13575_ (.CLK(clknet_leaf_86_clk),
    .D(_00121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[26] ));
 sky130_fd_sc_hd__dfxtp_4 _13576_ (.CLK(clknet_leaf_86_clk),
    .D(_00122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13577_ (.CLK(clknet_leaf_81_clk),
    .D(_00123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13578_ (.CLK(clknet_leaf_78_clk),
    .D(_00124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13579_ (.CLK(clknet_leaf_78_clk),
    .D(_00125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[30] ));
 sky130_fd_sc_hd__dfxtp_4 _13580_ (.CLK(clknet_leaf_78_clk),
    .D(_00126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.a_in[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13581_ (.CLK(clknet_leaf_74_clk),
    .D(_00127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13582_ (.CLK(clknet_leaf_73_clk),
    .D(_00128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13583_ (.CLK(clknet_leaf_73_clk),
    .D(_00129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13584_ (.CLK(clknet_leaf_51_clk),
    .D(_00130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13585_ (.CLK(clknet_leaf_51_clk),
    .D(_00131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13586_ (.CLK(clknet_leaf_59_clk),
    .D(_00132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13587_ (.CLK(clknet_leaf_59_clk),
    .D(_00133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13588_ (.CLK(clknet_leaf_59_clk),
    .D(_00134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13589_ (.CLK(clknet_leaf_61_clk),
    .D(_00135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13590_ (.CLK(clknet_leaf_63_clk),
    .D(_00136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13591_ (.CLK(clknet_leaf_63_clk),
    .D(_00137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13592_ (.CLK(clknet_leaf_63_clk),
    .D(_00138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13593_ (.CLK(clknet_leaf_64_clk),
    .D(_00139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13594_ (.CLK(clknet_leaf_67_clk),
    .D(_00140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13595_ (.CLK(clknet_leaf_67_clk),
    .D(_00141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13596_ (.CLK(clknet_leaf_68_clk),
    .D(_00142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13597_ (.CLK(clknet_leaf_69_clk),
    .D(_00143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13598_ (.CLK(clknet_leaf_69_clk),
    .D(_00144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13599_ (.CLK(clknet_leaf_69_clk),
    .D(_00145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13600_ (.CLK(clknet_leaf_84_clk),
    .D(_00146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13601_ (.CLK(clknet_leaf_85_clk),
    .D(_00147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13602_ (.CLK(clknet_leaf_86_clk),
    .D(_00148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13603_ (.CLK(clknet_leaf_87_clk),
    .D(_00149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13604_ (.CLK(clknet_leaf_86_clk),
    .D(_00150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13605_ (.CLK(clknet_leaf_81_clk),
    .D(_00151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13606_ (.CLK(clknet_leaf_80_clk),
    .D(_00152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13607_ (.CLK(clknet_leaf_79_clk),
    .D(_00153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13608_ (.CLK(clknet_leaf_78_clk),
    .D(_00154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13609_ (.CLK(clknet_leaf_78_clk),
    .D(_00155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13610_ (.CLK(clknet_leaf_82_clk),
    .D(_00156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13611_ (.CLK(clknet_leaf_74_clk),
    .D(_00157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13612_ (.CLK(clknet_leaf_71_clk),
    .D(_00158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.b_in[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13613_ (.CLK(clknet_leaf_74_clk),
    .D(_00159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13614_ (.CLK(clknet_leaf_73_clk),
    .D(_00160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13615_ (.CLK(clknet_leaf_73_clk),
    .D(_00161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13616_ (.CLK(clknet_leaf_51_clk),
    .D(_00162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13617_ (.CLK(clknet_leaf_51_clk),
    .D(_00163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13618_ (.CLK(clknet_leaf_59_clk),
    .D(_00164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13619_ (.CLK(clknet_leaf_59_clk),
    .D(_00165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13620_ (.CLK(clknet_leaf_59_clk),
    .D(_00166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13621_ (.CLK(clknet_leaf_61_clk),
    .D(_00167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13622_ (.CLK(clknet_leaf_63_clk),
    .D(_00168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13623_ (.CLK(clknet_leaf_63_clk),
    .D(_00169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13624_ (.CLK(clknet_leaf_63_clk),
    .D(_00170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13625_ (.CLK(clknet_leaf_64_clk),
    .D(_00171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13626_ (.CLK(clknet_leaf_67_clk),
    .D(_00172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13627_ (.CLK(clknet_leaf_67_clk),
    .D(_00173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13628_ (.CLK(clknet_leaf_68_clk),
    .D(_00174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13629_ (.CLK(clknet_leaf_68_clk),
    .D(_00175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13630_ (.CLK(clknet_leaf_69_clk),
    .D(_00176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13631_ (.CLK(clknet_leaf_84_clk),
    .D(_00177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_leaf_84_clk),
    .D(_00178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_leaf_85_clk),
    .D(_00179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_leaf_86_clk),
    .D(_00180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_leaf_87_clk),
    .D(_00181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_leaf_86_clk),
    .D(_00182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_leaf_81_clk),
    .D(_00183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_leaf_80_clk),
    .D(_00184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_leaf_79_clk),
    .D(_00185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_leaf_78_clk),
    .D(_00186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_leaf_82_clk),
    .D(_00187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_leaf_82_clk),
    .D(_00188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_leaf_74_clk),
    .D(_00189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_leaf_71_clk),
    .D(_00190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.c_in[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_leaf_71_clk),
    .D(_00191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_leaf_74_clk),
    .D(_00192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_leaf_73_clk),
    .D(_00193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_leaf_51_clk),
    .D(_00194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_leaf_60_clk),
    .D(_00195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13650_ (.CLK(clknet_leaf_60_clk),
    .D(_00196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_leaf_59_clk),
    .D(_00197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_4_15_0_clk),
    .D(_00198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13653_ (.CLK(clknet_leaf_61_clk),
    .D(_00199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13654_ (.CLK(clknet_leaf_63_clk),
    .D(_00200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_leaf_63_clk),
    .D(_00201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_leaf_64_clk),
    .D(_00202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_leaf_64_clk),
    .D(_00203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13658_ (.CLK(clknet_leaf_67_clk),
    .D(_00204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_leaf_67_clk),
    .D(_00205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_leaf_68_clk),
    .D(_00206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_leaf_68_clk),
    .D(_00207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13662_ (.CLK(clknet_leaf_69_clk),
    .D(_00208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_leaf_84_clk),
    .D(_00209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_leaf_84_clk),
    .D(_00210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_leaf_85_clk),
    .D(_00211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_leaf_87_clk),
    .D(_00212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13667_ (.CLK(clknet_leaf_87_clk),
    .D(_00213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13668_ (.CLK(clknet_leaf_87_clk),
    .D(_00214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13669_ (.CLK(clknet_leaf_88_clk),
    .D(_00215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13670_ (.CLK(clknet_leaf_80_clk),
    .D(_00216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13671_ (.CLK(clknet_leaf_80_clk),
    .D(_00217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13672_ (.CLK(clknet_leaf_78_clk),
    .D(_00218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13673_ (.CLK(clknet_leaf_82_clk),
    .D(_00219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13674_ (.CLK(clknet_leaf_82_clk),
    .D(_00220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13675_ (.CLK(clknet_leaf_71_clk),
    .D(_00221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13676_ (.CLK(clknet_leaf_71_clk),
    .D(_00222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.d_in[31] ));
 sky130_fd_sc_hd__dfxtp_4 _13677_ (.CLK(clknet_leaf_72_clk),
    .D(_00223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[0] ));
 sky130_fd_sc_hd__dfxtp_4 _13678_ (.CLK(clknet_leaf_71_clk),
    .D(_00224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[1] ));
 sky130_fd_sc_hd__dfxtp_4 _13679_ (.CLK(clknet_leaf_72_clk),
    .D(_00225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[2] ));
 sky130_fd_sc_hd__dfxtp_4 _13680_ (.CLK(clknet_leaf_66_clk),
    .D(_00226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[3] ));
 sky130_fd_sc_hd__dfxtp_4 _13681_ (.CLK(clknet_leaf_66_clk),
    .D(_00227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[4] ));
 sky130_fd_sc_hd__dfxtp_4 _13682_ (.CLK(clknet_leaf_66_clk),
    .D(_00228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[5] ));
 sky130_fd_sc_hd__dfxtp_4 _13683_ (.CLK(clknet_leaf_65_clk),
    .D(_00229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[6] ));
 sky130_fd_sc_hd__dfxtp_4 _13684_ (.CLK(clknet_leaf_65_clk),
    .D(_00230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[7] ));
 sky130_fd_sc_hd__dfxtp_4 _13685_ (.CLK(clknet_leaf_65_clk),
    .D(_00231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[8] ));
 sky130_fd_sc_hd__dfxtp_4 _13686_ (.CLK(clknet_leaf_65_clk),
    .D(_00232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[9] ));
 sky130_fd_sc_hd__dfxtp_4 _13687_ (.CLK(clknet_leaf_65_clk),
    .D(_00233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13688_ (.CLK(clknet_leaf_65_clk),
    .D(_00234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13689_ (.CLK(clknet_leaf_64_clk),
    .D(_00235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13690_ (.CLK(clknet_leaf_64_clk),
    .D(_00236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[13] ));
 sky130_fd_sc_hd__dfxtp_4 _13691_ (.CLK(clknet_leaf_67_clk),
    .D(_00237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[14] ));
 sky130_fd_sc_hd__dfxtp_4 _13692_ (.CLK(clknet_leaf_67_clk),
    .D(_00238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[15] ));
 sky130_fd_sc_hd__dfxtp_4 _13693_ (.CLK(clknet_leaf_68_clk),
    .D(_00239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[16] ));
 sky130_fd_sc_hd__dfxtp_4 _13694_ (.CLK(clknet_leaf_67_clk),
    .D(_00240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[17] ));
 sky130_fd_sc_hd__dfxtp_4 _13695_ (.CLK(clknet_leaf_68_clk),
    .D(_00241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[18] ));
 sky130_fd_sc_hd__dfxtp_4 _13696_ (.CLK(clknet_leaf_68_clk),
    .D(_00242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[19] ));
 sky130_fd_sc_hd__dfxtp_4 _13697_ (.CLK(clknet_leaf_83_clk),
    .D(_00243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[20] ));
 sky130_fd_sc_hd__dfxtp_4 _13698_ (.CLK(clknet_leaf_84_clk),
    .D(_00244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[21] ));
 sky130_fd_sc_hd__dfxtp_4 _13699_ (.CLK(clknet_leaf_85_clk),
    .D(_00245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[22] ));
 sky130_fd_sc_hd__dfxtp_4 _13700_ (.CLK(clknet_leaf_85_clk),
    .D(_00246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[23] ));
 sky130_fd_sc_hd__dfxtp_4 _13701_ (.CLK(clknet_leaf_83_clk),
    .D(_00247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[24] ));
 sky130_fd_sc_hd__dfxtp_4 _13702_ (.CLK(clknet_leaf_83_clk),
    .D(_00248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[25] ));
 sky130_fd_sc_hd__dfxtp_4 _13703_ (.CLK(clknet_leaf_83_clk),
    .D(_00249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[26] ));
 sky130_fd_sc_hd__dfxtp_4 _13704_ (.CLK(clknet_leaf_83_clk),
    .D(_00250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[27] ));
 sky130_fd_sc_hd__dfxtp_4 _13705_ (.CLK(clknet_leaf_83_clk),
    .D(_00251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[28] ));
 sky130_fd_sc_hd__dfxtp_4 _13706_ (.CLK(clknet_leaf_82_clk),
    .D(_00252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[29] ));
 sky130_fd_sc_hd__dfxtp_4 _13707_ (.CLK(clknet_leaf_82_clk),
    .D(_00253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[30] ));
 sky130_fd_sc_hd__dfxtp_4 _13708_ (.CLK(clknet_leaf_82_clk),
    .D(_00254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.e_in[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_leaf_70_clk),
    .D(_00255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13710_ (.CLK(clknet_leaf_71_clk),
    .D(_00256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_leaf_73_clk),
    .D(_00257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_leaf_66_clk),
    .D(_00258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_leaf_65_clk),
    .D(_00259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_leaf_60_clk),
    .D(_00260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_leaf_61_clk),
    .D(_00261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_leaf_61_clk),
    .D(_00262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_leaf_65_clk),
    .D(_00263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_leaf_65_clk),
    .D(_00264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_leaf_65_clk),
    .D(_00265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13720_ (.CLK(clknet_leaf_65_clk),
    .D(_00266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_leaf_65_clk),
    .D(_00267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_leaf_67_clk),
    .D(_00268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_leaf_67_clk),
    .D(_00269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_leaf_68_clk),
    .D(_00270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_leaf_68_clk),
    .D(_00271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_leaf_70_clk),
    .D(_00272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_leaf_69_clk),
    .D(_00273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_leaf_84_clk),
    .D(_00274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13729_ (.CLK(clknet_leaf_83_clk),
    .D(_00275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13730_ (.CLK(clknet_leaf_83_clk),
    .D(_00276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13731_ (.CLK(clknet_leaf_83_clk),
    .D(_00277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13732_ (.CLK(clknet_leaf_83_clk),
    .D(_00278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13733_ (.CLK(clknet_leaf_83_clk),
    .D(_00279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_leaf_81_clk),
    .D(_00280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_leaf_83_clk),
    .D(_00281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_leaf_83_clk),
    .D(_00282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13737_ (.CLK(clknet_leaf_70_clk),
    .D(_00283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_leaf_83_clk),
    .D(_00284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13739_ (.CLK(clknet_leaf_70_clk),
    .D(_00285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13740_ (.CLK(clknet_leaf_70_clk),
    .D(_00286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.f_in[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13741_ (.CLK(clknet_leaf_70_clk),
    .D(_00287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13742_ (.CLK(clknet_leaf_71_clk),
    .D(_00288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13743_ (.CLK(clknet_leaf_73_clk),
    .D(_00289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13744_ (.CLK(clknet_leaf_66_clk),
    .D(_00290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13745_ (.CLK(clknet_leaf_66_clk),
    .D(_00291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13746_ (.CLK(clknet_leaf_60_clk),
    .D(_00292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13747_ (.CLK(clknet_leaf_60_clk),
    .D(_00293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13748_ (.CLK(clknet_leaf_61_clk),
    .D(_00294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13749_ (.CLK(clknet_leaf_65_clk),
    .D(_00295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13750_ (.CLK(clknet_leaf_65_clk),
    .D(_00296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13751_ (.CLK(clknet_leaf_63_clk),
    .D(_00297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13752_ (.CLK(clknet_leaf_65_clk),
    .D(_00298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13753_ (.CLK(clknet_leaf_64_clk),
    .D(_00299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13754_ (.CLK(clknet_leaf_67_clk),
    .D(_00300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13755_ (.CLK(clknet_leaf_67_clk),
    .D(_00301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13756_ (.CLK(clknet_leaf_68_clk),
    .D(_00302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13757_ (.CLK(clknet_leaf_68_clk),
    .D(_00303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13758_ (.CLK(clknet_leaf_70_clk),
    .D(_00304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13759_ (.CLK(clknet_leaf_69_clk),
    .D(_00305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13760_ (.CLK(clknet_leaf_84_clk),
    .D(_00306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13761_ (.CLK(clknet_leaf_84_clk),
    .D(_00307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13762_ (.CLK(clknet_leaf_84_clk),
    .D(_00308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13763_ (.CLK(clknet_leaf_84_clk),
    .D(_00309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13764_ (.CLK(clknet_leaf_85_clk),
    .D(_00310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13765_ (.CLK(clknet_leaf_81_clk),
    .D(_00311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13766_ (.CLK(clknet_leaf_81_clk),
    .D(_00312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13767_ (.CLK(clknet_leaf_82_clk),
    .D(_00313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13768_ (.CLK(clknet_leaf_83_clk),
    .D(_00314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13769_ (.CLK(clknet_leaf_82_clk),
    .D(_00315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13770_ (.CLK(clknet_leaf_82_clk),
    .D(_00316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13771_ (.CLK(clknet_leaf_71_clk),
    .D(_00317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13772_ (.CLK(clknet_leaf_70_clk),
    .D(_00318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.g_in[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13773_ (.CLK(clknet_leaf_70_clk),
    .D(_00319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13774_ (.CLK(clknet_leaf_71_clk),
    .D(_00320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13775_ (.CLK(clknet_leaf_73_clk),
    .D(_00321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13776_ (.CLK(clknet_leaf_66_clk),
    .D(_00322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13777_ (.CLK(clknet_leaf_66_clk),
    .D(_00323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13778_ (.CLK(clknet_leaf_60_clk),
    .D(_00324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13779_ (.CLK(clknet_leaf_60_clk),
    .D(_00325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13780_ (.CLK(clknet_leaf_61_clk),
    .D(_00326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13781_ (.CLK(clknet_leaf_65_clk),
    .D(_00327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13782_ (.CLK(clknet_leaf_64_clk),
    .D(_00328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13783_ (.CLK(clknet_leaf_63_clk),
    .D(_00329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13784_ (.CLK(clknet_leaf_63_clk),
    .D(_00330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13785_ (.CLK(clknet_leaf_64_clk),
    .D(_00331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13786_ (.CLK(clknet_leaf_67_clk),
    .D(_00332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13787_ (.CLK(clknet_leaf_67_clk),
    .D(_00333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13788_ (.CLK(clknet_leaf_68_clk),
    .D(_00334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13789_ (.CLK(clknet_leaf_68_clk),
    .D(_00335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13790_ (.CLK(clknet_leaf_69_clk),
    .D(_00336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13791_ (.CLK(clknet_leaf_69_clk),
    .D(_00337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13792_ (.CLK(clknet_leaf_84_clk),
    .D(_00338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13793_ (.CLK(clknet_leaf_84_clk),
    .D(_00339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13794_ (.CLK(clknet_leaf_85_clk),
    .D(_00340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13795_ (.CLK(clknet_leaf_85_clk),
    .D(_00341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13796_ (.CLK(clknet_leaf_85_clk),
    .D(_00342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13797_ (.CLK(clknet_leaf_88_clk),
    .D(_00343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13798_ (.CLK(clknet_leaf_81_clk),
    .D(_00344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13799_ (.CLK(clknet_leaf_83_clk),
    .D(_00345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_81_clk),
    .D(_00346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13801_ (.CLK(clknet_leaf_82_clk),
    .D(_00347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_82_clk),
    .D(_00348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13803_ (.CLK(clknet_leaf_70_clk),
    .D(_00349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13804_ (.CLK(clknet_leaf_70_clk),
    .D(_00350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_out_digest.h_in[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13805_ (.CLK(clknet_leaf_49_clk),
    .D(_00351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_48_clk),
    .D(_00352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_49_clk),
    .D(_00353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13808_ (.CLK(clknet_leaf_49_clk),
    .D(_00354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13809_ (.CLK(clknet_leaf_47_clk),
    .D(_00355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13810_ (.CLK(clknet_leaf_47_clk),
    .D(_00356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13811_ (.CLK(clknet_leaf_49_clk),
    .D(_00357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13812_ (.CLK(clknet_leaf_47_clk),
    .D(_00358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13813_ (.CLK(clknet_leaf_49_clk),
    .D(_00359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13814_ (.CLK(clknet_leaf_47_clk),
    .D(_00360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13815_ (.CLK(clknet_leaf_48_clk),
    .D(_00361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13816_ (.CLK(clknet_leaf_48_clk),
    .D(_00362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13817_ (.CLK(clknet_leaf_48_clk),
    .D(_00363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13818_ (.CLK(clknet_leaf_48_clk),
    .D(_00364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13819_ (.CLK(clknet_leaf_47_clk),
    .D(_00365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13820_ (.CLK(clknet_leaf_48_clk),
    .D(_00366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13821_ (.CLK(clknet_leaf_48_clk),
    .D(_00367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13822_ (.CLK(clknet_leaf_48_clk),
    .D(_00368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13823_ (.CLK(clknet_leaf_76_clk),
    .D(_00369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13824_ (.CLK(clknet_leaf_76_clk),
    .D(_00370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13825_ (.CLK(clknet_leaf_110_clk),
    .D(_00371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13826_ (.CLK(clknet_leaf_110_clk),
    .D(_00372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13827_ (.CLK(clknet_leaf_110_clk),
    .D(_00373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13828_ (.CLK(clknet_leaf_110_clk),
    .D(_00374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[23] ));
 sky130_fd_sc_hd__dfxtp_2 _13829_ (.CLK(clknet_leaf_109_clk),
    .D(_00375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13830_ (.CLK(clknet_leaf_76_clk),
    .D(_00376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[25] ));
 sky130_fd_sc_hd__dfxtp_2 _13831_ (.CLK(clknet_leaf_76_clk),
    .D(_00377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13832_ (.CLK(clknet_leaf_76_clk),
    .D(_00378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13833_ (.CLK(clknet_leaf_110_clk),
    .D(_00379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13834_ (.CLK(clknet_leaf_76_clk),
    .D(_00380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13835_ (.CLK(clknet_leaf_76_clk),
    .D(_00381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13836_ (.CLK(clknet_leaf_76_clk),
    .D(_00382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_14[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_18_clk),
    .D(_00383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_17_clk),
    .D(_00384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_18_clk),
    .D(_00385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_18_clk),
    .D(_00386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_18_clk),
    .D(_00387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_18_clk),
    .D(_00388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13843_ (.CLK(clknet_leaf_17_clk),
    .D(_00389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_17_clk),
    .D(_00390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_17_clk),
    .D(_00391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_17_clk),
    .D(_00392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_21_clk),
    .D(_00393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_21_clk),
    .D(_00394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_21_clk),
    .D(_00395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_17_clk),
    .D(_00396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_21_clk),
    .D(_00397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_21_clk),
    .D(_00398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_22_clk),
    .D(_00399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_17_clk),
    .D(_00400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_22_clk),
    .D(_00401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_22_clk),
    .D(_00402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_23_clk),
    .D(_00403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_23_clk),
    .D(_00404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_23_clk),
    .D(_00405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_23_clk),
    .D(_00406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_23_clk),
    .D(_00407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_23_clk),
    .D(_00408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_22_clk),
    .D(_00409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_22_clk),
    .D(_00410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_21_clk),
    .D(_00411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13866_ (.CLK(clknet_leaf_21_clk),
    .D(_00412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_21_clk),
    .D(_00413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_18_clk),
    .D(_00414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_13[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_20_clk),
    .D(_00415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13870_ (.CLK(clknet_leaf_20_clk),
    .D(_00416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_21_clk),
    .D(_00417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_18_clk),
    .D(_00418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_19_clk),
    .D(_00419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13874_ (.CLK(clknet_leaf_18_clk),
    .D(_00420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13875_ (.CLK(clknet_leaf_20_clk),
    .D(_00421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_20_clk),
    .D(_00422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_20_clk),
    .D(_00423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13878_ (.CLK(clknet_leaf_22_clk),
    .D(_00424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_20_clk),
    .D(_00425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_22_clk),
    .D(_00426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_23_clk),
    .D(_00427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_23_clk),
    .D(_00428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_24_clk),
    .D(_00429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_24_clk),
    .D(_00430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13885_ (.CLK(clknet_leaf_24_clk),
    .D(_00431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_24_clk),
    .D(_00432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_24_clk),
    .D(_00433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13888_ (.CLK(clknet_leaf_24_clk),
    .D(_00434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_24_clk),
    .D(_00435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_24_clk),
    .D(_00436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_24_clk),
    .D(_00437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_24_clk),
    .D(_00438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_24_clk),
    .D(_00439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_24_clk),
    .D(_00440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_22_clk),
    .D(_00441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_22_clk),
    .D(_00442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_23_clk),
    .D(_00443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_22_clk),
    .D(_00444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_20_clk),
    .D(_00445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_18_clk),
    .D(_00446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_12[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13901_ (.CLK(clknet_leaf_95_clk),
    .D(_00447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.counter_iteration[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_95_clk),
    .D(_00448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.counter_iteration[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13903_ (.CLK(clknet_leaf_96_clk),
    .D(_00449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.counter_iteration[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13904_ (.CLK(clknet_leaf_105_clk),
    .D(_00450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.counter_iteration[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13905_ (.CLK(clknet_leaf_105_clk),
    .D(_00451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.counter_iteration[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_96_clk),
    .D(_00452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.counter_iteration[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_97_clk),
    .D(_00453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.counter_iteration[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_96_clk),
    .D(_00454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.counter_iteration[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_96_clk),
    .D(_00455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.counter_iteration[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_96_clk),
    .D(_00456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.counter_iteration[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_95_clk),
    .D(_00457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.counter_iteration[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13912_ (.CLK(clknet_leaf_105_clk),
    .D(_00458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.counter_iteration[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_105_clk),
    .D(_00459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.temp_case ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_46_clk),
    .D(_00460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_45_clk),
    .D(_00461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_45_clk),
    .D(_00462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_45_clk),
    .D(_00463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_44_clk),
    .D(_00464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13919_ (.CLK(clknet_leaf_44_clk),
    .D(_00465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_44_clk),
    .D(_00466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_44_clk),
    .D(_00467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_44_clk),
    .D(_00468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13923_ (.CLK(clknet_leaf_44_clk),
    .D(_00469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13924_ (.CLK(clknet_leaf_44_clk),
    .D(_00470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13925_ (.CLK(clknet_leaf_43_clk),
    .D(_00471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13926_ (.CLK(clknet_leaf_44_clk),
    .D(_00472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13927_ (.CLK(clknet_leaf_43_clk),
    .D(_00473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13928_ (.CLK(clknet_leaf_53_clk),
    .D(_00474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13929_ (.CLK(clknet_leaf_52_clk),
    .D(_00475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_52_clk),
    .D(_00476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_52_clk),
    .D(_00477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13932_ (.CLK(clknet_leaf_52_clk),
    .D(_00478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_50_clk),
    .D(_00479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13934_ (.CLK(clknet_leaf_50_clk),
    .D(_00480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13935_ (.CLK(clknet_leaf_52_clk),
    .D(_00481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_53_clk),
    .D(_00482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_53_clk),
    .D(_00483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_50_clk),
    .D(_00484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_43_clk),
    .D(_00485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_49_clk),
    .D(_00486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_46_clk),
    .D(_00487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_46_clk),
    .D(_00488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_46_clk),
    .D(_00489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_43_clk),
    .D(_00490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_43_clk),
    .D(_00491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_43_clk),
    .D(_00492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_53_clk),
    .D(_00493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _13948_ (.CLK(clknet_leaf_53_clk),
    .D(_00494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _13949_ (.CLK(clknet_leaf_54_clk),
    .D(_00495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _13950_ (.CLK(clknet_leaf_54_clk),
    .D(_00496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13951_ (.CLK(clknet_leaf_54_clk),
    .D(_00497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13952_ (.CLK(clknet_leaf_54_clk),
    .D(_00498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13953_ (.CLK(clknet_leaf_52_clk),
    .D(_00499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13954_ (.CLK(clknet_leaf_54_clk),
    .D(_00500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13955_ (.CLK(clknet_leaf_52_clk),
    .D(_00501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13956_ (.CLK(clknet_leaf_52_clk),
    .D(_00502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13957_ (.CLK(clknet_leaf_59_clk),
    .D(_00503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _13958_ (.CLK(clknet_leaf_59_clk),
    .D(_00504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13959_ (.CLK(clknet_leaf_58_clk),
    .D(_00505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13960_ (.CLK(clknet_leaf_59_clk),
    .D(_00506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13961_ (.CLK(clknet_leaf_58_clk),
    .D(_00507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13962_ (.CLK(clknet_leaf_59_clk),
    .D(_00508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13963_ (.CLK(clknet_leaf_55_clk),
    .D(_00509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _13964_ (.CLK(clknet_leaf_55_clk),
    .D(_00510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13965_ (.CLK(clknet_leaf_57_clk),
    .D(_00511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _13966_ (.CLK(clknet_leaf_55_clk),
    .D(_00512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13967_ (.CLK(clknet_leaf_55_clk),
    .D(_00513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _13968_ (.CLK(clknet_leaf_54_clk),
    .D(_00514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _13969_ (.CLK(clknet_leaf_53_clk),
    .D(_00515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _13970_ (.CLK(clknet_leaf_54_clk),
    .D(_00516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _13971_ (.CLK(clknet_leaf_42_clk),
    .D(_00517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[25] ));
 sky130_fd_sc_hd__dfxtp_2 _13972_ (.CLK(clknet_leaf_42_clk),
    .D(_00518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[26] ));
 sky130_fd_sc_hd__dfxtp_2 _13973_ (.CLK(clknet_leaf_42_clk),
    .D(_00519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[27] ));
 sky130_fd_sc_hd__dfxtp_2 _13974_ (.CLK(clknet_leaf_42_clk),
    .D(_00520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _13975_ (.CLK(clknet_leaf_42_clk),
    .D(_00521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _13976_ (.CLK(clknet_leaf_42_clk),
    .D(_00522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _13977_ (.CLK(clknet_leaf_42_clk),
    .D(_00523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13978_ (.CLK(clknet_leaf_42_clk),
    .D(_00524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13979_ (.CLK(clknet_leaf_54_clk),
    .D(_00525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13980_ (.CLK(clknet_leaf_55_clk),
    .D(_00526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13981_ (.CLK(clknet_leaf_55_clk),
    .D(_00527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13982_ (.CLK(clknet_leaf_55_clk),
    .D(_00528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13983_ (.CLK(clknet_leaf_55_clk),
    .D(_00529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_56_clk),
    .D(_00530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_57_clk),
    .D(_00531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_56_clk),
    .D(_00532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13987_ (.CLK(clknet_leaf_57_clk),
    .D(_00533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13988_ (.CLK(clknet_leaf_57_clk),
    .D(_00534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13989_ (.CLK(clknet_leaf_58_clk),
    .D(_00535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13990_ (.CLK(clknet_leaf_57_clk),
    .D(_00536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13991_ (.CLK(clknet_leaf_58_clk),
    .D(_00537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13992_ (.CLK(clknet_leaf_58_clk),
    .D(_00538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13993_ (.CLK(clknet_leaf_57_clk),
    .D(_00539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13994_ (.CLK(clknet_leaf_58_clk),
    .D(_00540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13995_ (.CLK(clknet_leaf_57_clk),
    .D(_00541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13996_ (.CLK(clknet_leaf_57_clk),
    .D(_00542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13997_ (.CLK(clknet_leaf_56_clk),
    .D(_00543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13998_ (.CLK(clknet_leaf_56_clk),
    .D(_00544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13999_ (.CLK(clknet_leaf_56_clk),
    .D(_00545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14000_ (.CLK(clknet_leaf_56_clk),
    .D(_00546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14001_ (.CLK(clknet_leaf_55_clk),
    .D(_00547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14002_ (.CLK(clknet_leaf_40_clk),
    .D(_00548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14003_ (.CLK(clknet_leaf_41_clk),
    .D(_00549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14004_ (.CLK(clknet_leaf_40_clk),
    .D(_00550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14005_ (.CLK(clknet_leaf_41_clk),
    .D(_00551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14006_ (.CLK(clknet_leaf_41_clk),
    .D(_00552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14007_ (.CLK(clknet_leaf_41_clk),
    .D(_00553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14008_ (.CLK(clknet_leaf_41_clk),
    .D(_00554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14009_ (.CLK(clknet_leaf_42_clk),
    .D(_00555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14010_ (.CLK(clknet_leaf_42_clk),
    .D(_00556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14011_ (.CLK(clknet_leaf_42_clk),
    .D(_00557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14012_ (.CLK(clknet_leaf_41_clk),
    .D(_00558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14013_ (.CLK(clknet_leaf_41_clk),
    .D(_00559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14014_ (.CLK(clknet_leaf_41_clk),
    .D(_00560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14015_ (.CLK(clknet_leaf_56_clk),
    .D(_00561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14016_ (.CLK(clknet_leaf_40_clk),
    .D(_00562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14017_ (.CLK(clknet_leaf_40_clk),
    .D(_00563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14018_ (.CLK(clknet_leaf_56_clk),
    .D(_00564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14019_ (.CLK(clknet_leaf_56_clk),
    .D(_00565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14020_ (.CLK(clknet_leaf_56_clk),
    .D(_00566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14021_ (.CLK(clknet_leaf_57_clk),
    .D(_00567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14022_ (.CLK(clknet_leaf_56_clk),
    .D(_00568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14023_ (.CLK(clknet_leaf_57_clk),
    .D(_00569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14024_ (.CLK(clknet_leaf_57_clk),
    .D(_00570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14025_ (.CLK(clknet_leaf_56_clk),
    .D(_00571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14026_ (.CLK(clknet_leaf_56_clk),
    .D(_00572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14027_ (.CLK(clknet_leaf_56_clk),
    .D(_00573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14028_ (.CLK(clknet_leaf_56_clk),
    .D(_00574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14029_ (.CLK(clknet_leaf_56_clk),
    .D(_00575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14030_ (.CLK(clknet_leaf_40_clk),
    .D(_00576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14031_ (.CLK(clknet_leaf_40_clk),
    .D(_00577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14032_ (.CLK(clknet_leaf_40_clk),
    .D(_00578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14033_ (.CLK(clknet_leaf_40_clk),
    .D(_00579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14034_ (.CLK(clknet_leaf_40_clk),
    .D(_00580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14035_ (.CLK(clknet_leaf_39_clk),
    .D(_00581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14036_ (.CLK(clknet_leaf_39_clk),
    .D(_00582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14037_ (.CLK(clknet_leaf_39_clk),
    .D(_00583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14038_ (.CLK(clknet_leaf_39_clk),
    .D(_00584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14039_ (.CLK(clknet_leaf_41_clk),
    .D(_00585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14040_ (.CLK(clknet_leaf_41_clk),
    .D(_00586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14041_ (.CLK(clknet_leaf_44_clk),
    .D(_00587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_3[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14042_ (.CLK(clknet_leaf_44_clk),
    .D(_00588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14043_ (.CLK(clknet_leaf_42_clk),
    .D(_00589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14044_ (.CLK(clknet_leaf_42_clk),
    .D(_00590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14045_ (.CLK(clknet_leaf_41_clk),
    .D(_00591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14046_ (.CLK(clknet_leaf_39_clk),
    .D(_00592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14047_ (.CLK(clknet_leaf_39_clk),
    .D(_00593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14048_ (.CLK(clknet_leaf_39_clk),
    .D(_00594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14049_ (.CLK(clknet_leaf_40_clk),
    .D(_00595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14050_ (.CLK(clknet_leaf_39_clk),
    .D(_00596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14051_ (.CLK(clknet_leaf_40_clk),
    .D(_00597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14052_ (.CLK(clknet_leaf_40_clk),
    .D(_00598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14053_ (.CLK(clknet_leaf_40_clk),
    .D(_00599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14054_ (.CLK(clknet_leaf_40_clk),
    .D(_00600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14055_ (.CLK(clknet_leaf_39_clk),
    .D(_00601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14056_ (.CLK(clknet_leaf_40_clk),
    .D(_00602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14057_ (.CLK(clknet_leaf_40_clk),
    .D(_00603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14058_ (.CLK(clknet_leaf_39_clk),
    .D(_00604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14059_ (.CLK(clknet_leaf_39_clk),
    .D(_00605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14060_ (.CLK(clknet_leaf_39_clk),
    .D(_00606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14061_ (.CLK(clknet_leaf_38_clk),
    .D(_00607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14062_ (.CLK(clknet_leaf_38_clk),
    .D(_00608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14063_ (.CLK(clknet_leaf_39_clk),
    .D(_00609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14064_ (.CLK(clknet_leaf_38_clk),
    .D(_00610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14065_ (.CLK(clknet_leaf_39_clk),
    .D(_00611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14066_ (.CLK(clknet_leaf_38_clk),
    .D(_00612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14067_ (.CLK(clknet_leaf_38_clk),
    .D(_00613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14068_ (.CLK(clknet_leaf_38_clk),
    .D(_00614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14069_ (.CLK(clknet_leaf_36_clk),
    .D(_00615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14070_ (.CLK(clknet_leaf_38_clk),
    .D(_00616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14071_ (.CLK(clknet_leaf_36_clk),
    .D(_00617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14072_ (.CLK(clknet_leaf_36_clk),
    .D(_00618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14073_ (.CLK(clknet_leaf_44_clk),
    .D(_00619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_4[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14074_ (.CLK(clknet_leaf_44_clk),
    .D(_00620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14075_ (.CLK(clknet_leaf_44_clk),
    .D(_00621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14076_ (.CLK(clknet_leaf_36_clk),
    .D(_00622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14077_ (.CLK(clknet_leaf_36_clk),
    .D(_00623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14078_ (.CLK(clknet_leaf_36_clk),
    .D(_00624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14079_ (.CLK(clknet_leaf_36_clk),
    .D(_00625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14080_ (.CLK(clknet_leaf_36_clk),
    .D(_00626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14081_ (.CLK(clknet_leaf_37_clk),
    .D(_00627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14082_ (.CLK(clknet_leaf_38_clk),
    .D(_00628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14083_ (.CLK(clknet_leaf_37_clk),
    .D(_00629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14084_ (.CLK(clknet_leaf_37_clk),
    .D(_00630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14085_ (.CLK(clknet_leaf_37_clk),
    .D(_00631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14086_ (.CLK(clknet_leaf_37_clk),
    .D(_00632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14087_ (.CLK(clknet_leaf_38_clk),
    .D(_00633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14088_ (.CLK(clknet_leaf_37_clk),
    .D(_00634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14089_ (.CLK(clknet_leaf_37_clk),
    .D(_00635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14090_ (.CLK(clknet_leaf_33_clk),
    .D(_00636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14091_ (.CLK(clknet_leaf_37_clk),
    .D(_00637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14092_ (.CLK(clknet_leaf_37_clk),
    .D(_00638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14093_ (.CLK(clknet_leaf_32_clk),
    .D(_00639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14094_ (.CLK(clknet_leaf_32_clk),
    .D(_00640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14095_ (.CLK(clknet_leaf_33_clk),
    .D(_00641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14096_ (.CLK(clknet_leaf_33_clk),
    .D(_00642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14097_ (.CLK(clknet_leaf_33_clk),
    .D(_00643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14098_ (.CLK(clknet_leaf_33_clk),
    .D(_00644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14099_ (.CLK(clknet_leaf_36_clk),
    .D(_00645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14100_ (.CLK(clknet_leaf_37_clk),
    .D(_00646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14101_ (.CLK(clknet_leaf_33_clk),
    .D(_00647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14102_ (.CLK(clknet_leaf_33_clk),
    .D(_00648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14103_ (.CLK(clknet_leaf_35_clk),
    .D(_00649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14104_ (.CLK(clknet_leaf_36_clk),
    .D(_00650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14105_ (.CLK(clknet_leaf_35_clk),
    .D(_00651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_5[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14106_ (.CLK(clknet_leaf_36_clk),
    .D(_00652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14107_ (.CLK(clknet_leaf_36_clk),
    .D(_00653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14108_ (.CLK(clknet_leaf_36_clk),
    .D(_00654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14109_ (.CLK(clknet_leaf_36_clk),
    .D(_00655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14110_ (.CLK(clknet_leaf_36_clk),
    .D(_00656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14111_ (.CLK(clknet_leaf_36_clk),
    .D(_00657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14112_ (.CLK(clknet_leaf_36_clk),
    .D(_00658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14113_ (.CLK(clknet_leaf_37_clk),
    .D(_00659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14114_ (.CLK(clknet_leaf_37_clk),
    .D(_00660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14115_ (.CLK(clknet_leaf_37_clk),
    .D(_00661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14116_ (.CLK(clknet_leaf_37_clk),
    .D(_00662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14117_ (.CLK(clknet_leaf_37_clk),
    .D(_00663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14118_ (.CLK(clknet_leaf_32_clk),
    .D(_00664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14119_ (.CLK(clknet_leaf_32_clk),
    .D(_00665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14120_ (.CLK(clknet_leaf_32_clk),
    .D(_00666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14121_ (.CLK(clknet_leaf_32_clk),
    .D(_00667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14122_ (.CLK(clknet_leaf_32_clk),
    .D(_00668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14123_ (.CLK(clknet_leaf_32_clk),
    .D(_00669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14124_ (.CLK(clknet_leaf_32_clk),
    .D(_00670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_32_clk),
    .D(_00671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_32_clk),
    .D(_00672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14127_ (.CLK(clknet_leaf_32_clk),
    .D(_00673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_33_clk),
    .D(_00674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_34_clk),
    .D(_00675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_34_clk),
    .D(_00676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_33_clk),
    .D(_00677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_34_clk),
    .D(_00678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_34_clk),
    .D(_00679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_34_clk),
    .D(_00680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_34_clk),
    .D(_00681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_34_clk),
    .D(_00682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_34_clk),
    .D(_00683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_6[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_35_clk),
    .D(_00684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_44_clk),
    .D(_00685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_36_clk),
    .D(_00686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_44_clk),
    .D(_00687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14142_ (.CLK(clknet_leaf_36_clk),
    .D(_00688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14143_ (.CLK(clknet_leaf_35_clk),
    .D(_00689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14144_ (.CLK(clknet_leaf_35_clk),
    .D(_00690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14145_ (.CLK(clknet_leaf_35_clk),
    .D(_00691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14146_ (.CLK(clknet_leaf_35_clk),
    .D(_00692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_35_clk),
    .D(_00693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_33_clk),
    .D(_00694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14149_ (.CLK(clknet_leaf_33_clk),
    .D(_00695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14150_ (.CLK(clknet_leaf_34_clk),
    .D(_00696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_31_clk),
    .D(_00697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_32_clk),
    .D(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_31_clk),
    .D(_00699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_31_clk),
    .D(_00700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_31_clk),
    .D(_00701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_32_clk),
    .D(_00702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_32_clk),
    .D(_00703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_31_clk),
    .D(_00704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_31_clk),
    .D(_00705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_31_clk),
    .D(_00706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_34_clk),
    .D(_00707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_34_clk),
    .D(_00708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_34_clk),
    .D(_00709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_34_clk),
    .D(_00710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_34_clk),
    .D(_00711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_34_clk),
    .D(_00712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_34_clk),
    .D(_00713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_34_clk),
    .D(_00714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_35_clk),
    .D(_00715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_7[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_35_clk),
    .D(_00716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_45_clk),
    .D(_00717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_45_clk),
    .D(_00718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_45_clk),
    .D(_00719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_45_clk),
    .D(_00720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_35_clk),
    .D(_00721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_35_clk),
    .D(_00722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_35_clk),
    .D(_00723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_35_clk),
    .D(_00724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_35_clk),
    .D(_00725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_35_clk),
    .D(_00726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_28_clk),
    .D(_00727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_28_clk),
    .D(_00728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_29_clk),
    .D(_00729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_29_clk),
    .D(_00730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_29_clk),
    .D(_00731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_29_clk),
    .D(_00732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_29_clk),
    .D(_00733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_29_clk),
    .D(_00734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_29_clk),
    .D(_00735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_29_clk),
    .D(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_31_clk),
    .D(_00737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_29_clk),
    .D(_00738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14193_ (.CLK(clknet_leaf_29_clk),
    .D(_00739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14194_ (.CLK(clknet_leaf_29_clk),
    .D(_00740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14195_ (.CLK(clknet_leaf_29_clk),
    .D(_00741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_29_clk),
    .D(_00742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_29_clk),
    .D(_00743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_28_clk),
    .D(_00744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_28_clk),
    .D(_00745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_28_clk),
    .D(_00746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_28_clk),
    .D(_00747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_8[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14202_ (.CLK(clknet_leaf_19_clk),
    .D(_00748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_45_clk),
    .D(_00749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14204_ (.CLK(clknet_leaf_45_clk),
    .D(_00750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_45_clk),
    .D(_00751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14206_ (.CLK(clknet_leaf_45_clk),
    .D(_00752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_45_clk),
    .D(_00753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14208_ (.CLK(clknet_leaf_28_clk),
    .D(_00754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_28_clk),
    .D(_00755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14210_ (.CLK(clknet_leaf_28_clk),
    .D(_00756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14211_ (.CLK(clknet_leaf_28_clk),
    .D(_00757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14212_ (.CLK(clknet_leaf_28_clk),
    .D(_00758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_28_clk),
    .D(_00759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_27_clk),
    .D(_00760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14215_ (.CLK(clknet_leaf_28_clk),
    .D(_00761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14216_ (.CLK(clknet_leaf_28_clk),
    .D(_00762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14217_ (.CLK(clknet_leaf_28_clk),
    .D(_00763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14218_ (.CLK(clknet_leaf_30_clk),
    .D(_00764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14219_ (.CLK(clknet_leaf_30_clk),
    .D(_00765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14220_ (.CLK(clknet_leaf_30_clk),
    .D(_00766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[18] ));
 sky130_fd_sc_hd__dfxtp_2 _14221_ (.CLK(clknet_leaf_30_clk),
    .D(_00767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[19] ));
 sky130_fd_sc_hd__dfxtp_2 _14222_ (.CLK(clknet_leaf_26_clk),
    .D(_00768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[20] ));
 sky130_fd_sc_hd__dfxtp_2 _14223_ (.CLK(clknet_leaf_26_clk),
    .D(_00769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[21] ));
 sky130_fd_sc_hd__dfxtp_2 _14224_ (.CLK(clknet_leaf_26_clk),
    .D(_00770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[22] ));
 sky130_fd_sc_hd__dfxtp_2 _14225_ (.CLK(clknet_leaf_26_clk),
    .D(_00771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[23] ));
 sky130_fd_sc_hd__dfxtp_2 _14226_ (.CLK(clknet_leaf_26_clk),
    .D(_00772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_26_clk),
    .D(_00773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[25] ));
 sky130_fd_sc_hd__dfxtp_2 _14228_ (.CLK(clknet_leaf_26_clk),
    .D(_00774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[26] ));
 sky130_fd_sc_hd__dfxtp_2 _14229_ (.CLK(clknet_leaf_27_clk),
    .D(_00775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_27_clk),
    .D(_00776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_27_clk),
    .D(_00777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_27_clk),
    .D(_00778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_19_clk),
    .D(_00779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_9[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_19_clk),
    .D(_00780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_19_clk),
    .D(_00781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_19_clk),
    .D(_00782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_19_clk),
    .D(_00783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_19_clk),
    .D(_00784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_19_clk),
    .D(_00785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_19_clk),
    .D(_00786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_19_clk),
    .D(_00787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_28_clk),
    .D(_00788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_28_clk),
    .D(_00789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_28_clk),
    .D(_00790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_27_clk),
    .D(_00791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_27_clk),
    .D(_00792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_26_clk),
    .D(_00793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_26_clk),
    .D(_00794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_26_clk),
    .D(_00795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_25_clk),
    .D(_00796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_25_clk),
    .D(_00797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_26_clk),
    .D(_00798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_25_clk),
    .D(_00799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_25_clk),
    .D(_00800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_26_clk),
    .D(_00801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_26_clk),
    .D(_00802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_25_clk),
    .D(_00803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_25_clk),
    .D(_00804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_26_clk),
    .D(_00805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_26_clk),
    .D(_00806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_27_clk),
    .D(_00807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_27_clk),
    .D(_00808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_20_clk),
    .D(_00809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_27_clk),
    .D(_00810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_20_clk),
    .D(_00811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_10[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_19_clk),
    .D(_00812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_19_clk),
    .D(_00813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_19_clk),
    .D(_00814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_18_clk),
    .D(_00815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_19_clk),
    .D(_00816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_19_clk),
    .D(_00817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_20_clk),
    .D(_00818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_20_clk),
    .D(_00819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_20_clk),
    .D(_00820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_20_clk),
    .D(_00821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_20_clk),
    .D(_00822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_27_clk),
    .D(_00823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_23_clk),
    .D(_00824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_23_clk),
    .D(_00825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_25_clk),
    .D(_00826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_25_clk),
    .D(_00827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_24_clk),
    .D(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_25_clk),
    .D(_00829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_24_clk),
    .D(_00830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_24_clk),
    .D(_00831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_24_clk),
    .D(_00832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_25_clk),
    .D(_00833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_25_clk),
    .D(_00834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_25_clk),
    .D(_00835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_25_clk),
    .D(_00836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_25_clk),
    .D(_00837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_25_clk),
    .D(_00838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_27_clk),
    .D(_00839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_25_clk),
    .D(_00840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_20_clk),
    .D(_00841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_20_clk),
    .D(_00842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_20_clk),
    .D(_00843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.mreg_11[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_90_clk),
    .D(_00000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00036_));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_97_clk),
    .D(_00011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00047_));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_95_clk),
    .D(_00022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00058_));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_90_clk),
    .D(_00025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00061_));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_4_5_0_clk),
    .D(_00026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00062_));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_95_clk),
    .D(_00027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00063_));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_90_clk),
    .D(_00028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00064_));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_95_clk),
    .D(_00029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00065_));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_95_clk),
    .D(_00030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00066_));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_90_clk),
    .D(_00031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00067_));
 sky130_fd_sc_hd__dfxtp_1 _14308_ (.CLK(clknet_leaf_90_clk),
    .D(_00001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00037_));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_92_clk),
    .D(_00002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00038_));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_92_clk),
    .D(_00003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00039_));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_93_clk),
    .D(_00004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00040_));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.CLK(clknet_leaf_92_clk),
    .D(_00005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00041_));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_91_clk),
    .D(_00006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00042_));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_92_clk),
    .D(_00007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00043_));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_91_clk),
    .D(_00008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00044_));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.CLK(clknet_leaf_92_clk),
    .D(_00009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00045_));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_95_clk),
    .D(_00010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00046_));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_93_clk),
    .D(_00012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00048_));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.CLK(clknet_leaf_91_clk),
    .D(_00013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00049_));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.CLK(clknet_leaf_90_clk),
    .D(_00014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00050_));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_89_clk),
    .D(_00015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00051_));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_90_clk),
    .D(_00016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00052_));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_95_clk),
    .D(_00017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00053_));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_90_clk),
    .D(_00018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00054_));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_90_clk),
    .D(_00019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00055_));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_95_clk),
    .D(_00020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00056_));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_89_clk),
    .D(_00021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00057_));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_90_clk),
    .D(_00023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00059_));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_90_clk),
    .D(_00024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(_00060_));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_10_clk),
    .D(_00844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.m_size[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_114_clk),
    .D(_00845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.m_size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_2_clk),
    .D(_00846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.m_size[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_2_clk),
    .D(_00847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.m_size[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_124_clk),
    .D(_00848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.m_size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_10_clk),
    .D(_00849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.m_size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_10_clk),
    .D(_00850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.m_size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_105_clk),
    .D(_00851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.counter_iteration[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14338_ (.CLK(clknet_leaf_105_clk),
    .D(_00852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.msg_scheduler.counter_iteration[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14339_ (.CLK(clknet_leaf_111_clk),
    .D(_00853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14340_ (.CLK(clknet_leaf_111_clk),
    .D(_00854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_111_clk),
    .D(_00855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_111_clk),
    .D(_00856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14343_ (.CLK(clknet_leaf_112_clk),
    .D(_00857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out3[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14344_ (.CLK(clknet_leaf_112_clk),
    .D(_00858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out3[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14345_ (.CLK(clknet_leaf_111_clk),
    .D(_00859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_112_clk),
    .D(_00860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_108_clk),
    .D(_00861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_out3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_108_clk),
    .D(_00862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.flag_0_15 ));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.CLK(clknet_leaf_110_clk),
    .D(_00863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.CLK(clknet_leaf_9_clk),
    .D(_00864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.CLK(clknet_leaf_7_clk),
    .D(_00865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.CLK(clknet_leaf_14_clk),
    .D(_00866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_110_clk),
    .D(_00867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.CLK(clknet_leaf_14_clk),
    .D(_00868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.CLK(clknet_leaf_14_clk),
    .D(_00869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.CLK(clknet_leaf_11_clk),
    .D(_00870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_110_clk),
    .D(_00871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_110_clk),
    .D(_00872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_14_clk),
    .D(_00873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.CLK(clknet_leaf_14_clk),
    .D(_00874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.CLK(clknet_leaf_14_clk),
    .D(_00875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_14_clk),
    .D(_00876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_15_clk),
    .D(_00877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.CLK(clknet_leaf_109_clk),
    .D(_00878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_77_clk),
    .D(_00879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.CLK(clknet_leaf_77_clk),
    .D(_00880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.CLK(clknet_leaf_77_clk),
    .D(_00881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.CLK(clknet_leaf_77_clk),
    .D(_00882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.CLK(clknet_leaf_77_clk),
    .D(_00883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.CLK(clknet_leaf_109_clk),
    .D(_00884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14371_ (.CLK(clknet_leaf_77_clk),
    .D(_00885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14372_ (.CLK(clknet_leaf_110_clk),
    .D(_00886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_109_clk),
    .D(_00887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_110_clk),
    .D(_00888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_109_clk),
    .D(_00889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14376_ (.CLK(clknet_leaf_110_clk),
    .D(_00890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14377_ (.CLK(clknet_leaf_110_clk),
    .D(_00891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14378_ (.CLK(clknet_leaf_110_clk),
    .D(_00892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14379_ (.CLK(clknet_leaf_110_clk),
    .D(_00893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.CLK(clknet_leaf_110_clk),
    .D(_00894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.data_in_padd[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14381_ (.CLK(clknet_leaf_79_clk),
    .D(_00895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.hashing_done ));
 sky130_fd_sc_hd__dfxtp_4 _14382_ (.CLK(clknet_leaf_108_clk),
    .D(_00896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.padding_done ));
 sky130_fd_sc_hd__dfxtp_1 _14383_ (.CLK(clknet_leaf_107_clk),
    .D(_00897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.temp_chk ));
 sky130_fd_sc_hd__dfxtp_2 _14384_ (.CLK(clknet_leaf_47_clk),
    .D(_00898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14385_ (.CLK(clknet_leaf_47_clk),
    .D(_00899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14386_ (.CLK(clknet_leaf_47_clk),
    .D(_00900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14387_ (.CLK(clknet_leaf_47_clk),
    .D(_00901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14388_ (.CLK(clknet_leaf_47_clk),
    .D(_00902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14389_ (.CLK(clknet_leaf_15_clk),
    .D(_00903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[5] ));
 sky130_fd_sc_hd__dfxtp_4 _14390_ (.CLK(clknet_leaf_15_clk),
    .D(_00904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[6] ));
 sky130_fd_sc_hd__dfxtp_4 _14391_ (.CLK(clknet_leaf_15_clk),
    .D(_00905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[7] ));
 sky130_fd_sc_hd__dfxtp_4 _14392_ (.CLK(clknet_leaf_47_clk),
    .D(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[8] ));
 sky130_fd_sc_hd__dfxtp_4 _14393_ (.CLK(clknet_leaf_47_clk),
    .D(_00907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[9] ));
 sky130_fd_sc_hd__dfxtp_4 _14394_ (.CLK(clknet_leaf_47_clk),
    .D(_00908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[10] ));
 sky130_fd_sc_hd__dfxtp_4 _14395_ (.CLK(clknet_leaf_15_clk),
    .D(_00909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[11] ));
 sky130_fd_sc_hd__dfxtp_4 _14396_ (.CLK(clknet_leaf_47_clk),
    .D(_00910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[12] ));
 sky130_fd_sc_hd__dfxtp_4 _14397_ (.CLK(clknet_leaf_48_clk),
    .D(_00911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[13] ));
 sky130_fd_sc_hd__dfxtp_4 _14398_ (.CLK(clknet_leaf_47_clk),
    .D(_00912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[14] ));
 sky130_fd_sc_hd__dfxtp_4 _14399_ (.CLK(clknet_leaf_75_clk),
    .D(_00913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14400_ (.CLK(clknet_leaf_75_clk),
    .D(_00914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14401_ (.CLK(clknet_leaf_75_clk),
    .D(_00915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14402_ (.CLK(clknet_leaf_75_clk),
    .D(_00916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[18] ));
 sky130_fd_sc_hd__dfxtp_2 _14403_ (.CLK(clknet_leaf_76_clk),
    .D(_00917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[19] ));
 sky130_fd_sc_hd__dfxtp_4 _14404_ (.CLK(clknet_leaf_76_clk),
    .D(_00918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[20] ));
 sky130_fd_sc_hd__dfxtp_2 _14405_ (.CLK(clknet_leaf_76_clk),
    .D(_00919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[21] ));
 sky130_fd_sc_hd__dfxtp_2 _14406_ (.CLK(clknet_leaf_77_clk),
    .D(_00920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[22] ));
 sky130_fd_sc_hd__dfxtp_2 _14407_ (.CLK(clknet_leaf_77_clk),
    .D(_00921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[23] ));
 sky130_fd_sc_hd__dfxtp_2 _14408_ (.CLK(clknet_leaf_109_clk),
    .D(_00922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[24] ));
 sky130_fd_sc_hd__dfxtp_2 _14409_ (.CLK(clknet_leaf_77_clk),
    .D(_00923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[25] ));
 sky130_fd_sc_hd__dfxtp_2 _14410_ (.CLK(clknet_leaf_109_clk),
    .D(_00924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[26] ));
 sky130_fd_sc_hd__dfxtp_2 _14411_ (.CLK(clknet_leaf_109_clk),
    .D(_00925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[27] ));
 sky130_fd_sc_hd__dfxtp_2 _14412_ (.CLK(clknet_leaf_110_clk),
    .D(_00926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[28] ));
 sky130_fd_sc_hd__dfxtp_2 _14413_ (.CLK(clknet_leaf_110_clk),
    .D(_00927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[29] ));
 sky130_fd_sc_hd__dfxtp_2 _14414_ (.CLK(clknet_leaf_110_clk),
    .D(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_15_clk),
    .D(_00929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.iter_processing.w[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_107_clk),
    .D(_00930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_512_block[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14417_ (.CLK(clknet_leaf_107_clk),
    .D(_00931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_512_block[1] ));
 sky130_fd_sc_hd__dfxtp_4 _14418_ (.CLK(clknet_leaf_106_clk),
    .D(_00932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_512_block[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14419_ (.CLK(clknet_leaf_107_clk),
    .D(_00933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_512_block[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14420_ (.CLK(clknet_leaf_108_clk),
    .D(_00934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_512_block[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14421_ (.CLK(clknet_leaf_112_clk),
    .D(_00935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_512_block[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14422_ (.CLK(clknet_leaf_108_clk),
    .D(_00936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.add_512_block[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_120_clk),
    .D(_00937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_117_clk),
    .D(_00938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_100_clk),
    .D(_00939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.CLK(clknet_leaf_118_clk),
    .D(_00940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.CLK(clknet_leaf_100_clk),
    .D(_00941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.CLK(clknet_leaf_117_clk),
    .D(_00942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.CLK(clknet_leaf_119_clk),
    .D(_00943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14430_ (.CLK(clknet_leaf_116_clk),
    .D(_00944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.CLK(clknet_leaf_97_clk),
    .D(_00945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.CLK(clknet_leaf_96_clk),
    .D(_00946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_103_clk),
    .D(_00947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.CLK(clknet_leaf_104_clk),
    .D(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_96_clk),
    .D(_00949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.CLK(clknet_leaf_97_clk),
    .D(_00950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_97_clk),
    .D(_00951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_103_clk),
    .D(_00952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_8_clk),
    .D(_00953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.CLK(clknet_leaf_9_clk),
    .D(_00954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_11_clk),
    .D(_00955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_9_clk),
    .D(_00956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_9_clk),
    .D(_00957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_11_clk),
    .D(_00958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14445_ (.CLK(clknet_leaf_8_clk),
    .D(_00959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.CLK(clknet_leaf_112_clk),
    .D(_00960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_3_clk),
    .D(_00961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_9_clk),
    .D(_00962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_7_clk),
    .D(_00963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_6_clk),
    .D(_00964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.CLK(clknet_leaf_6_clk),
    .D(_00965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.CLK(clknet_leaf_5_clk),
    .D(_00966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.CLK(clknet_leaf_4_clk),
    .D(_00967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_112_clk),
    .D(_00968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_120_clk),
    .D(_00969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_119_clk),
    .D(_00970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_126_clk),
    .D(_00971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_126_clk),
    .D(_00972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_126_clk),
    .D(_00973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_126_clk),
    .D(_00974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_121_clk),
    .D(_00975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_115_clk),
    .D(_00976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_98_clk),
    .D(_00977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_98_clk),
    .D(_00978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_99_clk),
    .D(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_101_clk),
    .D(_00980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_98_clk),
    .D(_00981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_100_clk),
    .D(_00982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_98_clk),
    .D(_00983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_102_clk),
    .D(_00984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_13_clk),
    .D(_00985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_12_clk),
    .D(_00986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_12_clk),
    .D(_00987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_12_clk),
    .D(_00988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_9_clk),
    .D(_00989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_8_clk),
    .D(_00990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_8_clk),
    .D(_00991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_113_clk),
    .D(_00992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_6_clk),
    .D(_00993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_9_clk),
    .D(_00994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_7_clk),
    .D(_00995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_6_clk),
    .D(_00996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_6_clk),
    .D(_00997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_5_clk),
    .D(_00998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_4_clk),
    .D(_00999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_114_clk),
    .D(_01000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_120_clk),
    .D(_01001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_120_clk),
    .D(_01002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.CLK(clknet_leaf_121_clk),
    .D(_01003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.CLK(clknet_leaf_121_clk),
    .D(_01004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.CLK(clknet_leaf_121_clk),
    .D(_01005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_122_clk),
    .D(_01006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_121_clk),
    .D(_01007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_123_clk),
    .D(_01008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_104_clk),
    .D(_01009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_105_clk),
    .D(_01010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_104_clk),
    .D(_01011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_105_clk),
    .D(_01012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_103_clk),
    .D(_01013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_103_clk),
    .D(_01014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_105_clk),
    .D(_01015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_107_clk),
    .D(_01016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_13_clk),
    .D(_01017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_8_clk),
    .D(_01018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_16_clk),
    .D(_01019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_16_clk),
    .D(_01020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_8_clk),
    .D(_01021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_12_clk),
    .D(_01022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_22_clk),
    .D(_01023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_109_clk),
    .D(_01024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_4_clk),
    .D(_01025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_2_clk),
    .D(_01026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_2_clk),
    .D(_01027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_4_clk),
    .D(_01028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_4_clk),
    .D(_01029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_4_clk),
    .D(_01030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_3_clk),
    .D(_01031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_114_clk),
    .D(_01032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_122_clk),
    .D(_01033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_120_clk),
    .D(_01034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_126_clk),
    .D(_01035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_126_clk),
    .D(_01036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_125_clk),
    .D(_01037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_126_clk),
    .D(_01038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_121_clk),
    .D(_01039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_114_clk),
    .D(_01040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_79_clk),
    .D(_01041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_106_clk),
    .D(_01042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_106_clk),
    .D(_01043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_105_clk),
    .D(_01044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_106_clk),
    .D(_01045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.CLK(clknet_leaf_106_clk),
    .D(_01046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_106_clk),
    .D(_01047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_102_clk),
    .D(_01048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_8_clk),
    .D(_01049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_12_clk),
    .D(_01050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_12_clk),
    .D(_01051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_8_clk),
    .D(_01052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_9_clk),
    .D(_01053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_11_clk),
    .D(_01054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_8_clk),
    .D(_01055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_111_clk),
    .D(_01056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_6_clk),
    .D(_01057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_6_clk),
    .D(_01058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_7_clk),
    .D(_01059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_3_clk),
    .D(_01060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_5_clk),
    .D(_01061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_6_clk),
    .D(_01062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_9_clk),
    .D(_01063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_111_clk),
    .D(_01064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_119_clk),
    .D(_01065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_119_clk),
    .D(_01066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_119_clk),
    .D(_01067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_118_clk),
    .D(_01068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_119_clk),
    .D(_01069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_120_clk),
    .D(_01070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_119_clk),
    .D(_01071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_117_clk),
    .D(_01072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_96_clk),
    .D(_01073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_96_clk),
    .D(_01074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_96_clk),
    .D(_01075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_96_clk),
    .D(_01076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_96_clk),
    .D(_01077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_96_clk),
    .D(_01078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_98_clk),
    .D(_01079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_116_clk),
    .D(_01080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_16_clk),
    .D(_01081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_14_clk),
    .D(_01082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_16_clk),
    .D(_01083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_16_clk),
    .D(_01084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_21_clk),
    .D(_01085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_22_clk),
    .D(_01086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_16_clk),
    .D(_01087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_112_clk),
    .D(_01088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_0_clk),
    .D(_01089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_2_clk),
    .D(_01090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_4_clk),
    .D(_01091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_4_clk),
    .D(_01092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_5_clk),
    .D(_01093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_4_clk),
    .D(_01094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_leaf_4_clk),
    .D(_01095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.CLK(clknet_leaf_113_clk),
    .D(_01096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_122_clk),
    .D(_01097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_120_clk),
    .D(_01098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_118_clk),
    .D(_01099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.CLK(clknet_leaf_118_clk),
    .D(_01100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_118_clk),
    .D(_01101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.CLK(clknet_leaf_117_clk),
    .D(_01102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_117_clk),
    .D(_01103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_117_clk),
    .D(_01104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_98_clk),
    .D(_01105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_98_clk),
    .D(_01106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_104_clk),
    .D(_01107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_101_clk),
    .D(_01108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_104_clk),
    .D(_01109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_101_clk),
    .D(_01110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.CLK(clknet_leaf_98_clk),
    .D(_01111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.CLK(clknet_leaf_102_clk),
    .D(_01112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_15_clk),
    .D(_01113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_14_clk),
    .D(_01114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.CLK(clknet_leaf_14_clk),
    .D(_01115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_14_clk),
    .D(_01116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_14_clk),
    .D(_01117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_14_clk),
    .D(_01118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_15_clk),
    .D(_01119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_110_clk),
    .D(_01120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.CLK(clknet_leaf_0_clk),
    .D(_01121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.CLK(clknet_leaf_2_clk),
    .D(_01122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_1_clk),
    .D(_01123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_5_clk),
    .D(_01124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_5_clk),
    .D(_01125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_5_clk),
    .D(_01126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.CLK(clknet_leaf_0_clk),
    .D(_01127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.CLK(clknet_leaf_113_clk),
    .D(_01128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_123_clk),
    .D(_01129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_120_clk),
    .D(_01130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_121_clk),
    .D(_01131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_121_clk),
    .D(_01132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_126_clk),
    .D(_01133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_122_clk),
    .D(_01134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_121_clk),
    .D(_01135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.CLK(clknet_leaf_115_clk),
    .D(_01136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_97_clk),
    .D(_01137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_98_clk),
    .D(_01138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_98_clk),
    .D(_01139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_96_clk),
    .D(_01140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_98_clk),
    .D(_01141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_97_clk),
    .D(_01142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_97_clk),
    .D(_01143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_116_clk),
    .D(_01144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.CLK(clknet_leaf_13_clk),
    .D(_01145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_12_clk),
    .D(_01146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_16_clk),
    .D(_01147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_16_clk),
    .D(_01148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_8_clk),
    .D(_01149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_21_clk),
    .D(_01150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_12_clk),
    .D(_01151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_108_clk),
    .D(_01152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_9_clk),
    .D(_01153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_2_clk),
    .D(_01154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.CLK(clknet_leaf_2_clk),
    .D(_01155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_10_clk),
    .D(_01156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_3_clk),
    .D(_01157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_3_clk),
    .D(_01158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.CLK(clknet_leaf_3_clk),
    .D(_01159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.CLK(clknet_leaf_113_clk),
    .D(_01160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_123_clk),
    .D(_01161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_122_clk),
    .D(_01162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_123_clk),
    .D(_01163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_123_clk),
    .D(_01164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_123_clk),
    .D(_01165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_122_clk),
    .D(_01166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_123_clk),
    .D(_01167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_115_clk),
    .D(_01168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_98_clk),
    .D(_01169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_96_clk),
    .D(_01170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_98_clk),
    .D(_01171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_96_clk),
    .D(_01172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_98_clk),
    .D(_01173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_98_clk),
    .D(_01174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_98_clk),
    .D(_01175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_116_clk),
    .D(_01176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_13_clk),
    .D(_01177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_13_clk),
    .D(_01178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_13_clk),
    .D(_01179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_12_clk),
    .D(_01180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_13_clk),
    .D(_01181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_14_clk),
    .D(_01182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_12_clk),
    .D(_01183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_110_clk),
    .D(_01184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_0_clk),
    .D(_01185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_2_clk),
    .D(_01186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_2_clk),
    .D(_01187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_1_clk),
    .D(_01188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_1_clk),
    .D(_01189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_124_clk),
    .D(_01190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_1_clk),
    .D(_01191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_114_clk),
    .D(_01192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_119_clk),
    .D(_01193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_119_clk),
    .D(_01194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_121_clk),
    .D(_01195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_120_clk),
    .D(_01196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_121_clk),
    .D(_01197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_122_clk),
    .D(_01198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_122_clk),
    .D(_01199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_115_clk),
    .D(_01200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_104_clk),
    .D(_01201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_104_clk),
    .D(_01202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_103_clk),
    .D(_01203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_105_clk),
    .D(_01204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_103_clk),
    .D(_01205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_103_clk),
    .D(_01206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.CLK(clknet_leaf_104_clk),
    .D(_01207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.CLK(clknet_leaf_116_clk),
    .D(_01208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_8_clk),
    .D(_01209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.CLK(clknet_leaf_7_clk),
    .D(_01210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_7_clk),
    .D(_01211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.CLK(clknet_leaf_22_clk),
    .D(_01212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_7_clk),
    .D(_01213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_7_clk),
    .D(_01214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_22_clk),
    .D(_01215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.CLK(clknet_leaf_111_clk),
    .D(_01216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_0_clk),
    .D(_01217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_0_clk),
    .D(_01218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_1_clk),
    .D(_01219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_5_clk),
    .D(_01220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_5_clk),
    .D(_01221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_5_clk),
    .D(_01222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_2_clk),
    .D(_01223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_114_clk),
    .D(_01224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[35][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_120_clk),
    .D(_01225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_125_clk),
    .D(_01226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_126_clk),
    .D(_01227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_126_clk),
    .D(_01228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_125_clk),
    .D(_01229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_122_clk),
    .D(_01230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.CLK(clknet_leaf_121_clk),
    .D(_01231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.CLK(clknet_leaf_123_clk),
    .D(_01232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_100_clk),
    .D(_01233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_99_clk),
    .D(_01234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_99_clk),
    .D(_01235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.CLK(clknet_leaf_101_clk),
    .D(_01236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_99_clk),
    .D(_01237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_100_clk),
    .D(_01238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_100_clk),
    .D(_01239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_116_clk),
    .D(_01240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_12_clk),
    .D(_01241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_7_clk),
    .D(_01242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14729_ (.CLK(clknet_leaf_7_clk),
    .D(_01243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.CLK(clknet_leaf_7_clk),
    .D(_01244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_8_clk),
    .D(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.CLK(clknet_leaf_7_clk),
    .D(_01246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_7_clk),
    .D(_01247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_11_clk),
    .D(_01248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[38][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.CLK(clknet_leaf_4_clk),
    .D(_01249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_4_clk),
    .D(_01250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.CLK(clknet_leaf_0_clk),
    .D(_01251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.CLK(clknet_leaf_9_clk),
    .D(_01252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_5_clk),
    .D(_01253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14740_ (.CLK(clknet_leaf_5_clk),
    .D(_01254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.CLK(clknet_leaf_3_clk),
    .D(_01255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.CLK(clknet_leaf_11_clk),
    .D(_01256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[39][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_120_clk),
    .D(_01257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.CLK(clknet_leaf_120_clk),
    .D(_01258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_126_clk),
    .D(_01259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_125_clk),
    .D(_01260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_125_clk),
    .D(_01261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14748_ (.CLK(clknet_leaf_126_clk),
    .D(_01262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.CLK(clknet_leaf_122_clk),
    .D(_01263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.CLK(clknet_leaf_123_clk),
    .D(_01264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14751_ (.CLK(clknet_leaf_106_clk),
    .D(_01265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14752_ (.CLK(clknet_leaf_106_clk),
    .D(_01266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14753_ (.CLK(clknet_leaf_106_clk),
    .D(_01267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14754_ (.CLK(clknet_leaf_103_clk),
    .D(_01268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14755_ (.CLK(clknet_leaf_103_clk),
    .D(_01269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14756_ (.CLK(clknet_leaf_106_clk),
    .D(_01270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14757_ (.CLK(clknet_leaf_105_clk),
    .D(_01271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14758_ (.CLK(clknet_leaf_102_clk),
    .D(_01272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14759_ (.CLK(clknet_leaf_8_clk),
    .D(_01273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14760_ (.CLK(clknet_leaf_12_clk),
    .D(_01274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.CLK(clknet_leaf_16_clk),
    .D(_01275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14762_ (.CLK(clknet_leaf_17_clk),
    .D(_01276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.CLK(clknet_leaf_11_clk),
    .D(_01277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.CLK(clknet_leaf_8_clk),
    .D(_01278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.CLK(clknet_leaf_16_clk),
    .D(_01279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.CLK(clknet_leaf_113_clk),
    .D(_01280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.CLK(clknet_leaf_3_clk),
    .D(_01281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_1_clk),
    .D(_01282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_2_clk),
    .D(_01283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_2_clk),
    .D(_01284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_3_clk),
    .D(_01285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_3_clk),
    .D(_01286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_3_clk),
    .D(_01287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_114_clk),
    .D(_01288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14775_ (.CLK(clknet_leaf_125_clk),
    .D(_01289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_122_clk),
    .D(_01290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.CLK(clknet_leaf_121_clk),
    .D(_01291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_121_clk),
    .D(_01292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_125_clk),
    .D(_01293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.CLK(clknet_leaf_126_clk),
    .D(_01294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_121_clk),
    .D(_01295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14782_ (.CLK(clknet_leaf_123_clk),
    .D(_01296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.CLK(clknet_leaf_106_clk),
    .D(_01297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_106_clk),
    .D(_01298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_108_clk),
    .D(_01299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_107_clk),
    .D(_01300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.CLK(clknet_leaf_107_clk),
    .D(_01301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.CLK(clknet_leaf_106_clk),
    .D(_01302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.CLK(clknet_leaf_106_clk),
    .D(_01303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_116_clk),
    .D(_01304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.CLK(clknet_leaf_11_clk),
    .D(_01305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.CLK(clknet_leaf_13_clk),
    .D(_01306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.CLK(clknet_leaf_13_clk),
    .D(_01307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.CLK(clknet_leaf_12_clk),
    .D(_01308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_13_clk),
    .D(_01309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.CLK(clknet_leaf_14_clk),
    .D(_01310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.CLK(clknet_leaf_11_clk),
    .D(_01311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.CLK(clknet_leaf_111_clk),
    .D(_01312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.CLK(clknet_leaf_0_clk),
    .D(_01313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_0_clk),
    .D(_01314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_1_clk),
    .D(_01315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.CLK(clknet_leaf_2_clk),
    .D(_01316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.CLK(clknet_leaf_1_clk),
    .D(_01317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_1_clk),
    .D(_01318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.CLK(clknet_leaf_4_clk),
    .D(_01319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14806_ (.CLK(clknet_leaf_114_clk),
    .D(_01320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.CLK(clknet_leaf_119_clk),
    .D(_01321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.CLK(clknet_leaf_119_clk),
    .D(_01322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14809_ (.CLK(clknet_leaf_117_clk),
    .D(_01323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14810_ (.CLK(clknet_leaf_118_clk),
    .D(_01324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.CLK(clknet_leaf_119_clk),
    .D(_01325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14812_ (.CLK(clknet_leaf_117_clk),
    .D(_01326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.CLK(clknet_leaf_119_clk),
    .D(_01327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14814_ (.CLK(clknet_leaf_117_clk),
    .D(_01328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14815_ (.CLK(clknet_leaf_98_clk),
    .D(_01329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.CLK(clknet_leaf_96_clk),
    .D(_01330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14817_ (.CLK(clknet_leaf_103_clk),
    .D(_01331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.CLK(clknet_leaf_104_clk),
    .D(_01332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.CLK(clknet_leaf_104_clk),
    .D(_01333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.CLK(clknet_leaf_101_clk),
    .D(_01334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_98_clk),
    .D(_01335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_102_clk),
    .D(_01336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_13_clk),
    .D(_01337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_9_clk),
    .D(_01338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_7_clk),
    .D(_01339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_22_clk),
    .D(_01340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_7_clk),
    .D(_01341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.CLK(clknet_leaf_7_clk),
    .D(_01342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.CLK(clknet_leaf_8_clk),
    .D(_01343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14830_ (.CLK(clknet_leaf_113_clk),
    .D(_01344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14831_ (.CLK(clknet_leaf_1_clk),
    .D(_01345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.CLK(clknet_leaf_4_clk),
    .D(_01346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.CLK(clknet_leaf_2_clk),
    .D(_01347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.CLK(clknet_leaf_2_clk),
    .D(_01348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14835_ (.CLK(clknet_leaf_0_clk),
    .D(_01349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.CLK(clknet_leaf_1_clk),
    .D(_01350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.CLK(clknet_leaf_4_clk),
    .D(_01351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_10_clk),
    .D(_01352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.CLK(clknet_leaf_119_clk),
    .D(_01353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_119_clk),
    .D(_01354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_118_clk),
    .D(_01355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_117_clk),
    .D(_01356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14843_ (.CLK(clknet_leaf_118_clk),
    .D(_01357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14844_ (.CLK(clknet_leaf_115_clk),
    .D(_01358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14845_ (.CLK(clknet_leaf_119_clk),
    .D(_01359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14846_ (.CLK(clknet_leaf_115_clk),
    .D(_01360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14847_ (.CLK(clknet_leaf_98_clk),
    .D(_01361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.CLK(clknet_leaf_99_clk),
    .D(_01362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.CLK(clknet_leaf_99_clk),
    .D(_01363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14850_ (.CLK(clknet_leaf_101_clk),
    .D(_01364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14851_ (.CLK(clknet_leaf_98_clk),
    .D(_01365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.CLK(clknet_leaf_100_clk),
    .D(_01366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14853_ (.CLK(clknet_leaf_99_clk),
    .D(_01367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14854_ (.CLK(clknet_leaf_102_clk),
    .D(_01368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14855_ (.CLK(clknet_leaf_11_clk),
    .D(_01369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.CLK(clknet_leaf_9_clk),
    .D(_01370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.CLK(clknet_leaf_7_clk),
    .D(_01371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.CLK(clknet_leaf_7_clk),
    .D(_01372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.CLK(clknet_leaf_7_clk),
    .D(_01373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_7_clk),
    .D(_01374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_11_clk),
    .D(_01375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_11_clk),
    .D(_01376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.CLK(clknet_leaf_1_clk),
    .D(_01377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.CLK(clknet_leaf_1_clk),
    .D(_01378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.CLK(clknet_leaf_1_clk),
    .D(_01379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.CLK(clknet_leaf_1_clk),
    .D(_01380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.CLK(clknet_leaf_1_clk),
    .D(_01381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_1_clk),
    .D(_01382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_124_clk),
    .D(_01383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_123_clk),
    .D(_01384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_124_clk),
    .D(_01385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_125_clk),
    .D(_01386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_125_clk),
    .D(_01387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_125_clk),
    .D(_01388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_125_clk),
    .D(_01389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.CLK(clknet_leaf_125_clk),
    .D(_01390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.CLK(clknet_leaf_125_clk),
    .D(_01391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.CLK(clknet_leaf_117_clk),
    .D(_01392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.CLK(clknet_leaf_100_clk),
    .D(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_99_clk),
    .D(_01394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_99_clk),
    .D(_01395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_101_clk),
    .D(_01396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_99_clk),
    .D(_01397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_100_clk),
    .D(_01398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_99_clk),
    .D(_01399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_117_clk),
    .D(_01400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_123_clk),
    .D(_01401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_9_clk),
    .D(_01402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_10_clk),
    .D(_01403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_9_clk),
    .D(_01404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_9_clk),
    .D(_01405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_9_clk),
    .D(_01406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_10_clk),
    .D(_01407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_9_clk),
    .D(_01408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_0_clk),
    .D(_01409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.CLK(clknet_leaf_0_clk),
    .D(_01410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_0_clk),
    .D(_01411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_1_clk),
    .D(_01412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.CLK(clknet_leaf_1_clk),
    .D(_01413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.CLK(clknet_leaf_1_clk),
    .D(_01414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_124_clk),
    .D(_01415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_123_clk),
    .D(_01416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14903_ (.CLK(clknet_leaf_124_clk),
    .D(_01417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.CLK(clknet_leaf_125_clk),
    .D(_01418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.CLK(clknet_leaf_124_clk),
    .D(_01419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.CLK(clknet_leaf_125_clk),
    .D(_01420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14907_ (.CLK(clknet_leaf_125_clk),
    .D(_01421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.CLK(clknet_leaf_123_clk),
    .D(_01422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14909_ (.CLK(clknet_leaf_124_clk),
    .D(_01423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.CLK(clknet_leaf_117_clk),
    .D(_01424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_100_clk),
    .D(_01425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_99_clk),
    .D(_01426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.CLK(clknet_leaf_99_clk),
    .D(_01427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_101_clk),
    .D(_01428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_99_clk),
    .D(_01429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_100_clk),
    .D(_01430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_99_clk),
    .D(_01431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_117_clk),
    .D(_01432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_2_clk),
    .D(_01433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_10_clk),
    .D(_01434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.CLK(clknet_leaf_11_clk),
    .D(_01435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.CLK(clknet_leaf_9_clk),
    .D(_01436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14923_ (.CLK(clknet_leaf_9_clk),
    .D(_01437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.CLK(clknet_leaf_10_clk),
    .D(_01438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.CLK(clknet_leaf_10_clk),
    .D(_01439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.CLK(clknet_leaf_10_clk),
    .D(_01440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.m_pad_pars.block_512[62][7] ));
 sky130_fd_sc_hd__dfxtp_2 _14927_ (.CLK(clknet_leaf_90_clk),
    .D(_01441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14928_ (.CLK(clknet_leaf_95_clk),
    .D(_01442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14929_ (.CLK(clknet_leaf_95_clk),
    .D(_01443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14930_ (.CLK(clknet_leaf_89_clk),
    .D(_01444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14931_ (.CLK(clknet_leaf_89_clk),
    .D(_01445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[4] ));
 sky130_fd_sc_hd__dfxtp_4 _14932_ (.CLK(clknet_leaf_95_clk),
    .D(_01446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[5] ));
 sky130_fd_sc_hd__dfxtp_4 _14933_ (.CLK(clknet_leaf_89_clk),
    .D(_01447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[6] ));
 sky130_fd_sc_hd__dfxtp_4 _14934_ (.CLK(clknet_leaf_89_clk),
    .D(_01448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[7] ));
 sky130_fd_sc_hd__dfxtp_4 _14935_ (.CLK(clknet_leaf_88_clk),
    .D(_01449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[8] ));
 sky130_fd_sc_hd__dfxtp_4 _14936_ (.CLK(clknet_leaf_91_clk),
    .D(_01450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[9] ));
 sky130_fd_sc_hd__dfxtp_4 _14937_ (.CLK(clknet_leaf_91_clk),
    .D(_01451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[10] ));
 sky130_fd_sc_hd__dfxtp_4 _14938_ (.CLK(clknet_leaf_91_clk),
    .D(_01452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[11] ));
 sky130_fd_sc_hd__dfxtp_4 _14939_ (.CLK(clknet_leaf_91_clk),
    .D(_01453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[12] ));
 sky130_fd_sc_hd__dfxtp_4 _14940_ (.CLK(clknet_leaf_91_clk),
    .D(_01454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[13] ));
 sky130_fd_sc_hd__dfxtp_4 _14941_ (.CLK(clknet_leaf_91_clk),
    .D(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[14] ));
 sky130_fd_sc_hd__dfxtp_4 _14942_ (.CLK(clknet_leaf_91_clk),
    .D(_01456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14943_ (.CLK(clknet_leaf_91_clk),
    .D(_01457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14944_ (.CLK(clknet_leaf_91_clk),
    .D(_01458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14945_ (.CLK(clknet_leaf_91_clk),
    .D(_01459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[18] ));
 sky130_fd_sc_hd__dfxtp_2 _14946_ (.CLK(clknet_leaf_91_clk),
    .D(_01460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[19] ));
 sky130_fd_sc_hd__dfxtp_2 _14947_ (.CLK(clknet_leaf_91_clk),
    .D(_01461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[20] ));
 sky130_fd_sc_hd__dfxtp_2 _14948_ (.CLK(clknet_leaf_91_clk),
    .D(_01462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.CLK(clknet_leaf_91_clk),
    .D(_01463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[22] ));
 sky130_fd_sc_hd__dfxtp_2 _14950_ (.CLK(clknet_leaf_89_clk),
    .D(_01464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[23] ));
 sky130_fd_sc_hd__dfxtp_2 _14951_ (.CLK(clknet_leaf_90_clk),
    .D(_01465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_89_clk),
    .D(_01466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.CLK(clknet_leaf_90_clk),
    .D(_01467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.CLK(clknet_leaf_89_clk),
    .D(_01468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[27] ));
 sky130_fd_sc_hd__dfxtp_2 _14955_ (.CLK(clknet_leaf_105_clk),
    .D(_01469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14956_ (.CLK(clknet_leaf_89_clk),
    .D(_01470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[29] ));
 sky130_fd_sc_hd__dfxtp_2 _14957_ (.CLK(clknet_leaf_89_clk),
    .D(_01471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[30] ));
 sky130_fd_sc_hd__dfxtp_2 _14958_ (.CLK(clknet_leaf_90_clk),
    .D(_01472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.K[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.CLK(clknet_leaf_95_clk),
    .D(_01473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\sha256cu.temp_case ));
 sky130_fd_sc_hd__conb_1 password_cracker_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net261));
 sky130_fd_sc_hd__conb_1 password_cracker_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net262));
 sky130_fd_sc_hd__conb_1 password_cracker_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net263));
 sky130_fd_sc_hd__conb_1 password_cracker_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net264));
 sky130_fd_sc_hd__conb_1 password_cracker_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net265));
 sky130_fd_sc_hd__conb_1 password_cracker_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net266));
 sky130_fd_sc_hd__conb_1 password_cracker_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net267));
 sky130_fd_sc_hd__conb_1 password_cracker_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net268));
 sky130_fd_sc_hd__conb_1 password_cracker_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net269));
 sky130_fd_sc_hd__conb_1 password_cracker_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net270));
 sky130_fd_sc_hd__conb_1 password_cracker_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net271));
 sky130_fd_sc_hd__conb_1 password_cracker_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net272));
 sky130_fd_sc_hd__conb_1 password_cracker_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net273));
 sky130_fd_sc_hd__conb_1 password_cracker_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net274));
 sky130_fd_sc_hd__conb_1 password_cracker_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net275));
 sky130_fd_sc_hd__conb_1 password_cracker_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net276));
 sky130_fd_sc_hd__conb_1 password_cracker_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net277));
 sky130_fd_sc_hd__conb_1 password_cracker_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net278));
 sky130_fd_sc_hd__conb_1 password_cracker_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net279));
 sky130_fd_sc_hd__conb_1 password_cracker_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net280));
 sky130_fd_sc_hd__conb_1 password_cracker_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net281));
 sky130_fd_sc_hd__conb_1 password_cracker_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net282));
 sky130_fd_sc_hd__conb_1 password_cracker_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net283));
 sky130_fd_sc_hd__conb_1 password_cracker_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net284));
 sky130_fd_sc_hd__conb_1 password_cracker_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net285));
 sky130_fd_sc_hd__conb_1 password_cracker_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net286));
 sky130_fd_sc_hd__conb_1 password_cracker_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net287));
 sky130_fd_sc_hd__conb_1 password_cracker_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net288));
 sky130_fd_sc_hd__conb_1 password_cracker_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net289));
 sky130_fd_sc_hd__conb_1 password_cracker_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net290));
 sky130_fd_sc_hd__conb_1 password_cracker_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net291));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(hash[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(hash[100]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(hash[101]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(hash[102]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(hash[103]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(hash[104]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(hash[105]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(hash[106]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(hash[107]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(hash[108]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(hash[109]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(hash[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(hash[110]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(hash[111]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(hash[112]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(hash[113]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(hash[114]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(hash[115]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(hash[116]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(hash[117]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(hash[118]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(hash[119]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(hash[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(hash[120]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(hash[121]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(hash[122]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(hash[123]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(hash[124]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(hash[125]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(hash[126]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(hash[127]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(hash[128]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(hash[129]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(hash[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(hash[130]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(hash[131]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(hash[132]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(hash[133]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(hash[134]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(hash[135]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(hash[136]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(hash[137]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(hash[138]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(hash[139]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(hash[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(hash[140]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(hash[141]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(hash[142]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(hash[143]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(hash[144]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(hash[145]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(hash[146]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(hash[147]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(hash[148]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(hash[149]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(hash[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(hash[150]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(hash[151]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(hash[152]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(hash[153]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(hash[154]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(hash[155]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(hash[156]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(hash[157]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(hash[158]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(hash[159]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(hash[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(hash[160]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(hash[161]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 input70 (.A(hash[162]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(hash[163]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(hash[164]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input73 (.A(hash[165]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(hash[166]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(hash[167]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(hash[168]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(hash[169]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(hash[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_2 input79 (.A(hash[170]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(hash[171]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(hash[172]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(hash[173]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__buf_2 input83 (.A(hash[174]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(hash[175]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(hash[176]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(hash[177]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(hash[178]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(hash[179]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(hash[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(hash[180]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(hash[181]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(hash[182]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(hash[183]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__buf_4 input94 (.A(hash[184]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 input95 (.A(hash[185]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(hash[186]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(hash[187]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(hash[188]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(hash[189]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(hash[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(hash[190]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(hash[191]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(hash[192]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__buf_2 input104 (.A(hash[193]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__buf_2 input105 (.A(hash[194]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(hash[195]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(hash[196]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(hash[197]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(hash[198]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input110 (.A(hash[199]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(hash[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 input112 (.A(hash[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__buf_4 input113 (.A(hash[200]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(hash[201]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(hash[202]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(hash[203]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 input117 (.A(hash[204]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 input118 (.A(hash[205]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(hash[206]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__buf_4 input120 (.A(hash[207]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(hash[208]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(hash[209]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(hash[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__buf_2 input124 (.A(hash[210]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(hash[211]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(hash[212]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(hash[213]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(hash[214]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(hash[215]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(hash[216]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__buf_4 input131 (.A(hash[217]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 input132 (.A(hash[218]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__buf_2 input133 (.A(hash[219]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(hash[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(hash[220]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 input136 (.A(hash[221]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(hash[222]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(hash[223]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(hash[224]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 input140 (.A(hash[225]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 input141 (.A(hash[226]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__buf_2 input142 (.A(hash[227]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 input143 (.A(hash[228]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(hash[229]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 input145 (.A(hash[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(hash[230]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(hash[231]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(hash[232]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(hash[233]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 input150 (.A(hash[234]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 input151 (.A(hash[235]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(hash[236]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 input153 (.A(hash[237]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(hash[238]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__buf_2 input155 (.A(hash[239]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(hash[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(hash[240]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(hash[241]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(hash[242]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(hash[243]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__buf_2 input161 (.A(hash[244]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(hash[245]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(hash[246]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(hash[247]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(hash[248]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 input166 (.A(hash[249]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(hash[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__buf_2 input168 (.A(hash[250]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(hash[251]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(hash[252]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 input171 (.A(hash[253]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(hash[254]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 input173 (.A(hash[255]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__buf_4 input174 (.A(hash[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlymetal6s2s_1 input175 (.A(hash[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(hash[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 input177 (.A(hash[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__dlymetal6s2s_1 input178 (.A(hash[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlymetal6s2s_1 input179 (.A(hash[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(hash[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__buf_2 input181 (.A(hash[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(hash[32]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 input183 (.A(hash[33]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__buf_2 input184 (.A(hash[34]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(hash[35]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(hash[36]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(hash[37]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(hash[38]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__buf_2 input189 (.A(hash[39]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 input190 (.A(hash[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(hash[40]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(hash[41]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(hash[42]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 input194 (.A(hash[43]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(hash[44]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(hash[45]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 input197 (.A(hash[46]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__buf_2 input198 (.A(hash[47]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__buf_4 input199 (.A(hash[48]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__buf_2 input200 (.A(hash[49]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__buf_2 input201 (.A(hash[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(hash[50]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(hash[51]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s2s_1 input204 (.A(hash[52]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(hash[53]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 input206 (.A(hash[54]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__dlymetal6s2s_1 input207 (.A(hash[55]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(hash[56]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 input209 (.A(hash[57]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 input210 (.A(hash[58]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 input211 (.A(hash[59]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(hash[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(hash[60]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(hash[61]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(hash[62]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__dlymetal6s2s_1 input216 (.A(hash[63]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 input217 (.A(hash[64]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(hash[65]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__buf_4 input219 (.A(hash[66]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input220 (.A(hash[67]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(hash[68]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 input222 (.A(hash[69]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(hash[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 input224 (.A(hash[70]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__dlymetal6s2s_1 input225 (.A(hash[71]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(hash[72]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 input227 (.A(hash[73]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(hash[74]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 input229 (.A(hash[75]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(hash[76]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 input231 (.A(hash[77]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__buf_4 input232 (.A(hash[78]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(hash[79]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 input234 (.A(hash[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__buf_2 input235 (.A(hash[80]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(hash[81]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__buf_2 input237 (.A(hash[82]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 input238 (.A(hash[83]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__buf_2 input239 (.A(hash[84]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input240 (.A(hash[85]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 input241 (.A(hash[86]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 input242 (.A(hash[87]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(hash[88]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__buf_2 input244 (.A(hash[89]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__buf_4 input245 (.A(hash[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(hash[90]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 input247 (.A(hash[91]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__dlymetal6s2s_1 input248 (.A(hash[92]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 input249 (.A(hash[93]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 input250 (.A(hash[94]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__buf_2 input251 (.A(hash[95]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__buf_2 input252 (.A(hash[96]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 input253 (.A(hash[97]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 input254 (.A(hash[98]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__buf_2 input255 (.A(hash[99]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__dlymetal6s2s_1 input256 (.A(hash[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 input257 (.A(reset),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(cracked));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(done));
 sky130_fd_sc_hd__conb_1 password_cracker_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net260));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_2_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_8_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_10_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_11_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_9_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_14_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_15_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_13_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_12_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_7_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_5_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_4_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_6_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_3_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_1_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_0_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_01479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_01479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_01494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_01494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_01513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_01513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_01521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_01526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_01551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_01551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_01554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_01554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_01554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_01554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_01975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_04881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_05342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\sha256cu.iter_processing.w[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\sha256cu.msg_scheduler.mreg_14[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\sha256cu.msg_scheduler.mreg_9[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net179),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(net219),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(net252),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(net254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(_01543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\sha256cu.iter_processing.w[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(_01558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(net185),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(net207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign password_count[0] = net260;
 assign password_count[10] = net270;
 assign password_count[11] = net271;
 assign password_count[12] = net272;
 assign password_count[13] = net273;
 assign password_count[14] = net274;
 assign password_count[15] = net275;
 assign password_count[16] = net276;
 assign password_count[17] = net277;
 assign password_count[18] = net278;
 assign password_count[19] = net279;
 assign password_count[1] = net261;
 assign password_count[20] = net280;
 assign password_count[21] = net281;
 assign password_count[22] = net282;
 assign password_count[23] = net283;
 assign password_count[24] = net284;
 assign password_count[25] = net285;
 assign password_count[26] = net286;
 assign password_count[27] = net287;
 assign password_count[28] = net288;
 assign password_count[29] = net289;
 assign password_count[2] = net262;
 assign password_count[30] = net290;
 assign password_count[31] = net291;
 assign password_count[3] = net263;
 assign password_count[4] = net264;
 assign password_count[5] = net265;
 assign password_count[6] = net266;
 assign password_count[7] = net267;
 assign password_count[8] = net268;
 assign password_count[9] = net269;
endmodule
