* NGSPICE file created from password_cracker.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt password_cracker VGND VPWR clk cracked done hash[0] hash[100] hash[101] hash[102]
+ hash[103] hash[104] hash[105] hash[106] hash[107] hash[108] hash[109] hash[10] hash[110]
+ hash[111] hash[112] hash[113] hash[114] hash[115] hash[116] hash[117] hash[118]
+ hash[119] hash[11] hash[120] hash[121] hash[122] hash[123] hash[124] hash[125] hash[126]
+ hash[127] hash[128] hash[129] hash[12] hash[130] hash[131] hash[132] hash[133] hash[134]
+ hash[135] hash[136] hash[137] hash[138] hash[139] hash[13] hash[140] hash[141] hash[142]
+ hash[143] hash[144] hash[145] hash[146] hash[147] hash[148] hash[149] hash[14] hash[150]
+ hash[151] hash[152] hash[153] hash[154] hash[155] hash[156] hash[157] hash[158]
+ hash[159] hash[15] hash[160] hash[161] hash[162] hash[163] hash[164] hash[165] hash[166]
+ hash[167] hash[168] hash[169] hash[16] hash[170] hash[171] hash[172] hash[173] hash[174]
+ hash[175] hash[176] hash[177] hash[178] hash[179] hash[17] hash[180] hash[181] hash[182]
+ hash[183] hash[184] hash[185] hash[186] hash[187] hash[188] hash[189] hash[18] hash[190]
+ hash[191] hash[192] hash[193] hash[194] hash[195] hash[196] hash[197] hash[198]
+ hash[199] hash[19] hash[1] hash[200] hash[201] hash[202] hash[203] hash[204] hash[205]
+ hash[206] hash[207] hash[208] hash[209] hash[20] hash[210] hash[211] hash[212] hash[213]
+ hash[214] hash[215] hash[216] hash[217] hash[218] hash[219] hash[21] hash[220] hash[221]
+ hash[222] hash[223] hash[224] hash[225] hash[226] hash[227] hash[228] hash[229]
+ hash[22] hash[230] hash[231] hash[232] hash[233] hash[234] hash[235] hash[236] hash[237]
+ hash[238] hash[239] hash[23] hash[240] hash[241] hash[242] hash[243] hash[244] hash[245]
+ hash[246] hash[247] hash[248] hash[249] hash[24] hash[250] hash[251] hash[252] hash[253]
+ hash[254] hash[255] hash[25] hash[26] hash[27] hash[28] hash[29] hash[2] hash[30]
+ hash[31] hash[32] hash[33] hash[34] hash[35] hash[36] hash[37] hash[38] hash[39]
+ hash[3] hash[40] hash[41] hash[42] hash[43] hash[44] hash[45] hash[46] hash[47]
+ hash[48] hash[49] hash[4] hash[50] hash[51] hash[52] hash[53] hash[54] hash[55]
+ hash[56] hash[57] hash[58] hash[59] hash[5] hash[60] hash[61] hash[62] hash[63]
+ hash[64] hash[65] hash[66] hash[67] hash[68] hash[69] hash[6] hash[70] hash[71]
+ hash[72] hash[73] hash[74] hash[75] hash[76] hash[77] hash[78] hash[79] hash[7]
+ hash[80] hash[81] hash[82] hash[83] hash[84] hash[85] hash[86] hash[87] hash[88]
+ hash[89] hash[8] hash[90] hash[91] hash[92] hash[93] hash[94] hash[95] hash[96]
+ hash[97] hash[98] hash[99] hash[9] init password_count[0] password_count[10] password_count[11]
+ password_count[12] password_count[13] password_count[14] password_count[15] password_count[16]
+ password_count[17] password_count[18] password_count[19] password_count[1] password_count[20]
+ password_count[21] password_count[22] password_count[23] password_count[24] password_count[25]
+ password_count[26] password_count[27] password_count[28] password_count[29] password_count[2]
+ password_count[30] password_count[31] password_count[3] password_count[4] password_count[5]
+ password_count[6] password_count[7] password_count[8] password_count[9] reset
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09671_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__buf_2
XFILLER_67_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06883_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__buf_6
XFILLER_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08622_ sha256cu.m_out_digest.c_in\[6\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[6\]
+ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__o22a_1
X_08553_ _03117_ _03119_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__and2b_1
X_07504_ sha256cu.m_out_digest.h_in\[3\] _02130_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08484_ sha256cu.m_out_digest.h_in\[28\] _03042_ _03084_ VGND VGND VPWR VPWR _03085_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07435_ _02005_ _02015_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__nor2_4
XFILLER_149_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07366_ _01986_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__buf_4
XFILLER_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09105_ _03588_ _03589_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__and2_1
X_07297_ sha256cu.m_pad_pars.add_512_block\[1\] _01939_ VGND VGND VPWR VPWR _01941_
+ sky130_fd_sc_hd__or2_2
X_09036_ _03489_ _03505_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__and3_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09938_ sha256cu.msg_scheduler.mreg_1\[8\] _04174_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__or2_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09869_ sha256cu.msg_scheduler.mreg_13\[20\] _04147_ VGND VGND VPWR VPWR _04159_
+ sky130_fd_sc_hd__or2_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _05718_ _05719_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__nor2_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12880_ sha256cu.m_pad_pars.block_512\[31\]\[0\] _06425_ VGND VGND VPWR VPWR _06426_
+ sky130_fd_sc_hd__and2_1
XANTENNA_213 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _05651_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__nand2_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_224 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_246 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14550_ clknet_leaf_111_clk _01064_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_268 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_235 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _05586_ _05566_ _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__a21oi_1
XANTENNA_279 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13501_ _01975_ _06764_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__and2_1
X_11693_ _05492_ _05507_ _05520_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__nand3_1
X_10713_ sha256cu.msg_scheduler.mreg_11\[21\] _04640_ VGND VGND VPWR VPWR _04643_
+ sky130_fd_sc_hd__or2_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ clknet_leaf_7_clk _00995_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10644_ sha256cu.msg_scheduler.mreg_10\[23\] _04601_ VGND VGND VPWR VPWR _04604_
+ sky130_fd_sc_hd__or2_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13432_ _06721_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10575_ sha256cu.msg_scheduler.mreg_8\[25\] _04554_ _04564_ _04557_ VGND VGND VPWR
+ VPWR _00741_ sky130_fd_sc_hd__o211a_1
X_13363_ _01923_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__buf_2
X_12314_ _05448_ _06115_ _06116_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__o21ai_1
XFILLER_108_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13294_ _06646_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12245_ sha256cu.data_in_padd\[27\] _05447_ _04053_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__a21o_1
XFILLER_5_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12176_ _05967_ _05984_ _05432_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11127_ sha256cu.m_pad_pars.block_512\[46\]\[0\] _04977_ _04981_ sha256cu.m_pad_pars.block_512\[54\]\[0\]
+ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__a221o_1
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11058_ _04808_ _04794_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__nor2_1
X_10009_ _04133_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14817_ clknet_leaf_103_clk _01331_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14748_ clknet_leaf_126_clk _01262_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14679_ clknet_leaf_119_clk _01193_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_07220_ _01584_ _01796_ _01872_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__or3_1
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07151_ _01679_ _01817_ _01818_ _01822_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__a31o_1
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07082_ _01602_ _01609_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__nor2_1
XFILLER_114_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07984_ sha256cu.m_out_digest.e_in\[22\] sha256cu.m_out_digest.e_in\[9\] VGND VGND
+ VPWR VPWR _02598_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09723_ sha256cu.msg_scheduler.mreg_14\[21\] _04073_ _04075_ _04064_ VGND VGND VPWR
+ VPWR _00372_ sky130_fd_sc_hd__o211a_1
X_06935_ _01625_ _01612_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__nand2_2
X_09654_ sha256cu.m_out_digest.h_in\[18\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[18\]
+ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__a22o_1
X_06866_ state\[1\] _01561_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__nand2_1
XFILLER_28_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08605_ sha256cu.m_out_digest.b_in\[23\] _03179_ _03178_ sha256cu.m_out_digest.a_in\[23\]
+ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__a22o_1
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09585_ sha256cu.m_out_digest.f_in\[25\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[25\]
+ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__o22a_1
X_06797_ net221 net225 net224 net227 VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__or4_2
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08536_ sha256cu.iter_processing.w\[29\] _03090_ _03135_ VGND VGND VPWR VPWR _03136_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_144_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08467_ _03035_ _03036_ _03067_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__or3b_1
XFILLER_23_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07418_ _02043_ _02044_ _02045_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__a21o_1
X_08398_ sha256cu.m_out_digest.e_in\[20\] _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__xnor2_4
XFILLER_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07349_ sha256cu.m_pad_pars.add_out0\[2\] _01961_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__and2_1
XFILLER_137_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10360_ sha256cu.msg_scheduler.mreg_6\[29\] _04441_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__or2_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10291_ sha256cu.msg_scheduler.mreg_4\[31\] _04393_ _04402_ _04397_ VGND VGND VPWR
+ VPWR _00619_ sky130_fd_sc_hd__o211a_1
XFILLER_128_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09019_ sha256cu.m_out_digest.h_in\[13\] sha256cu.m_out_digest.d_in\[13\] VGND VGND
+ VPWR VPWR _03508_ sky130_fd_sc_hd__and2_1
XFILLER_105_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12030_ sha256cu.iter_processing.w\[18\] _05666_ _05844_ _05640_ VGND VGND VPWR VPWR
+ _00916_ sky130_fd_sc_hd__o211a_1
XFILLER_132_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13981_ clknet_leaf_55_clk _00527_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12932_ sha256cu.m_pad_pars.block_512\[34\]\[0\] _06453_ VGND VGND VPWR VPWR _06454_
+ sky130_fd_sc_hd__and2_1
XFILLER_19_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ clknet_leaf_14_clk _01116_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12863_ sha256cu.m_pad_pars.block_512\[30\]\[0\] _06416_ VGND VGND VPWR VPWR _06417_
+ sky130_fd_sc_hd__and2_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _05636_ _05637_ _05465_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__a21oi_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12794_ _06251_ _05081_ _04961_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__or3_2
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ sha256cu.msg_scheduler.mreg_9\[7\] sha256cu.msg_scheduler.mreg_0\[7\] VGND
+ VGND VPWR VPWR _05571_ sky130_fd_sc_hd__nand2_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ clknet_leaf_106_clk _01047_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14464_ clknet_leaf_98_clk _00978_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11676_ sha256cu.iter_processing.w\[3\] _05430_ _05505_ _05335_ VGND VGND VPWR VPWR
+ _00901_ sky130_fd_sc_hd__o211a_1
X_13415_ sha256cu.m_pad_pars.block_512\[62\]\[4\] _01928_ VGND VGND VPWR VPWR _06709_
+ sky130_fd_sc_hd__and2_1
XFILLER_139_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10627_ _04580_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__buf_2
X_14395_ clknet_leaf_15_clk _00909_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[11\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_143_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10558_ sha256cu.msg_scheduler.mreg_9\[18\] _04548_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__or2_1
X_13346_ _06673_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13277_ _06637_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10489_ sha256cu.msg_scheduler.mreg_8\[21\] _04507_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__or2_1
X_12228_ sha256cu.msg_scheduler.mreg_9\[27\] sha256cu.msg_scheduler.mreg_0\[27\] VGND
+ VGND VPWR VPWR _06034_ sky130_fd_sc_hd__nand2_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12159_ sha256cu.msg_scheduler.mreg_9\[24\] sha256cu.msg_scheduler.mreg_0\[24\] VGND
+ VGND VPWR VPWR _05968_ sky130_fd_sc_hd__or2_1
XFILLER_69_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09370_ _02895_ _03813_ _03814_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__a21boi_1
X_08321_ _02900_ _02905_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand2_1
X_08252_ sha256cu.m_out_digest.g_in\[23\] sha256cu.m_out_digest.f_in\[23\] sha256cu.m_out_digest.e_in\[23\]
+ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__mux2_2
XFILLER_32_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07203_ _01823_ _01866_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__nand2_1
XFILLER_20_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_08183_ _02772_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07134_ _01666_ _01706_ _01646_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07065_ _01648_ _01687_ _01666_ _01745_ _01585_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__a311o_1
XFILLER_134_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07967_ sha256cu.K\[15\] _02581_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__xnor2_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09706_ sha256cu.iter_processing.w\[14\] _04054_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__or2_1
X_06918_ _01606_ _01609_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__nand2_2
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07898_ _02017_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__buf_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09637_ sha256cu.m_out_digest.h_in\[3\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[3\]
+ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__o22a_1
X_06849_ net2 net5 net4 net7 VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__or4_2
XFILLER_16_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09568_ sha256cu.m_out_digest.f_in\[10\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[10\]
+ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__a22o_1
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08519_ sha256cu.m_out_digest.e_in\[23\] _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__xnor2_4
XFILLER_70_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09499_ _03970_ _03971_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__nor2_1
X_11530_ sha256cu.m_pad_pars.block_512\[4\]\[5\] _05313_ _05299_ sha256cu.m_pad_pars.block_512\[12\]\[5\]
+ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__a22o_1
XFILLER_128_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11461_ _05293_ _05297_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__and3_2
XFILLER_152_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10412_ sha256cu.msg_scheduler.mreg_6\[19\] _04461_ _04471_ _04464_ VGND VGND VPWR
+ VPWR _00671_ sky130_fd_sc_hd__o211a_1
X_14180_ clknet_leaf_35_clk _00726_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13200_ _06596_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_1
X_11392_ _04747_ _05154_ _05155_ sha256cu.m_pad_pars.block_512\[21\]\[7\] VGND VGND
+ VPWR VPWR _05236_ sky130_fd_sc_hd__o22a_1
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10343_ sha256cu.msg_scheduler.mreg_6\[22\] _04428_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__or2_1
XFILLER_124_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13131_ _06559_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10274_ sha256cu.msg_scheduler.mreg_5\[25\] _04387_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__or2_1
X_13062_ _06522_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12013_ _05826_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__or2_1
XFILLER_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13964_ clknet_leaf_55_clk _00510_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_13895_ clknet_leaf_22_clk _00441_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12915_ sha256cu.m_pad_pars.block_512\[33\]\[0\] _06444_ VGND VGND VPWR VPWR _06445_
+ sky130_fd_sc_hd__and2_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12846_ sha256cu.m_pad_pars.block_512\[29\]\[0\] _06407_ VGND VGND VPWR VPWR _06408_
+ sky130_fd_sc_hd__and2_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ clknet_leaf_4_clk _01030_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12777_ _06251_ _05081_ _05130_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__or3_2
X_11728_ _05552_ _05554_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__xor2_1
XFILLER_119_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11659_ sha256cu.msg_scheduler.mreg_1\[21\] _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__xnor2_2
X_14447_ clknet_leaf_3_clk _00961_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14378_ clknet_leaf_110_clk _00892_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13329_ _06664_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08870_ sha256cu.m_out_digest.e_in\[7\] _02440_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__or2_1
XFILLER_85_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07821_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__buf_4
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07752_ sha256cu.m_out_digest.b_in\[10\] sha256cu.m_out_digest.a_in\[10\] VGND VGND
+ VPWR VPWR _02372_ sky130_fd_sc_hd__or2_1
XFILLER_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07683_ sha256cu.m_out_digest.a_in\[21\] sha256cu.m_out_digest.a_in\[10\] VGND VGND
+ VPWR VPWR _02305_ sky130_fd_sc_hd__xnor2_2
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09422_ _02113_ _03894_ _03897_ _02332_ sha256cu.m_out_digest.e_in\[26\] VGND VGND
+ VPWR VPWR _00249_ sky130_fd_sc_hd__a32o_1
X_09353_ _03804_ _03805_ _03802_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__a21o_1
XFILLER_61_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08304_ _02858_ _02859_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__and2b_1
XFILLER_33_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09284_ _03762_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__or2_1
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08235_ _02767_ _02840_ _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__o21ba_1
XFILLER_121_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08166_ sha256cu.m_out_digest.h_in\[21\] _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07117_ _01792_ _01653_ _01626_ _01659_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__o22a_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08097_ sha256cu.m_out_digest.g_in\[19\] sha256cu.m_out_digest.f_in\[19\] sha256cu.m_out_digest.e_in\[19\]
+ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__mux2_2
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07048_ _01730_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__inv_2
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08999_ _03475_ _03462_ _03488_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__o21ai_1
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10961_ _04756_ _04767_ _04827_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__and3_2
X_13680_ clknet_leaf_66_clk _00226_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_44_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12700_ sha256cu.m_pad_pars.block_512\[20\]\[4\] _06325_ VGND VGND VPWR VPWR _06330_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10892_ _04704_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__or2_2
X_12631_ _06293_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12562_ _06256_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12493_ sha256cu.m_pad_pars.block_512\[8\]\[4\] _06214_ VGND VGND VPWR VPWR _06219_
+ sky130_fd_sc_hd__and2_1
X_11513_ sha256cu.m_pad_pars.block_512\[52\]\[3\] _05310_ _05288_ sha256cu.m_pad_pars.block_512\[48\]\[3\]
+ _05352_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__a221o_1
X_14301_ clknet_leaf_90_clk _00025_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__dfxtp_1
X_14232_ clknet_leaf_27_clk _00778_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11444_ sha256cu.m_pad_pars.add_out0\[5\] sha256cu.m_pad_pars.add_out0\[4\] _01935_
+ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__and3_1
XFILLER_50_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14163_ clknet_leaf_34_clk _00709_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11375_ sha256cu.data_in_padd\[21\] _04741_ _04742_ _05220_ VGND VGND VPWR VPWR _00884_
+ sky130_fd_sc_hd__a22o_1
X_14094_ clknet_leaf_32_clk _00640_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10326_ sha256cu.msg_scheduler.mreg_5\[14\] _04421_ _04422_ _04410_ VGND VGND VPWR
+ VPWR _00634_ sky130_fd_sc_hd__o211a_1
X_13114_ _06550_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__clkbuf_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _04263_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__buf_2
XFILLER_112_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13045_ _06513_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__clkbuf_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10188_ _04263_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__buf_2
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13947_ clknet_leaf_53_clk _00493_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13878_ clknet_leaf_22_clk _00424_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12829_ sha256cu.m_pad_pars.block_512\[28\]\[0\] _06398_ VGND VGND VPWR VPWR _06399_
+ sky130_fd_sc_hd__and2_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08020_ _02610_ _02608_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__or2b_1
XFILLER_128_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ sha256cu.msg_scheduler.mreg_0\[22\] _04208_ _04219_ _04211_ VGND VGND VPWR
+ VPWR _00482_ sky130_fd_sc_hd__o211a_1
XFILLER_143_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08922_ _03413_ _03414_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__nor2_1
XFILLER_130_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08853_ sha256cu.K\[7\] _03347_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__xor2_1
XFILLER_112_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07804_ sha256cu.m_out_digest.h_in\[10\] _02384_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__nand2_1
X_08784_ _03280_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand2_1
XFILLER_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07735_ _02353_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07666_ sha256cu.K\[7\] _02288_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__xnor2_2
X_09405_ sha256cu.K\[26\] _03880_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__xnor2_1
X_07597_ sha256cu.iter_processing.w\[5\] _02192_ _02191_ VGND VGND VPWR VPWR _02221_
+ sky130_fd_sc_hd__a21o_1
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09336_ sha256cu.m_out_digest.h_in\[24\] sha256cu.m_out_digest.d_in\[24\] VGND VGND
+ VPWR VPWR _03814_ sky130_fd_sc_hd__nand2_1
X_09267_ _03746_ _03747_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__xnor2_1
X_08218_ _02782_ _02787_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__a21boi_1
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09198_ _03676_ _03680_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__nor2_1
XFILLER_5_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08149_ _02703_ _02725_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__nor2_1
X_11160_ sha256cu.data_in_padd\[8\] _04741_ _04742_ _05018_ VGND VGND VPWR VPWR _00871_
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10111_ sha256cu.msg_scheduler.mreg_2\[18\] _04288_ _04299_ _04291_ VGND VGND VPWR
+ VPWR _00542_ sky130_fd_sc_hd__o211a_1
XFILLER_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11091_ sha256cu.data_in_padd\[7\] _04840_ _04931_ _04950_ _01974_ VGND VGND VPWR
+ VPWR _00870_ sky130_fd_sc_hd__o221a_1
X_10042_ sha256cu.msg_scheduler.mreg_1\[21\] _04247_ _04259_ _04250_ VGND VGND VPWR
+ VPWR _00513_ sky130_fd_sc_hd__o211a_1
XFILLER_49_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14850_ clknet_leaf_101_clk _01364_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13801_ clknet_leaf_82_clk _00347_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14781_ clknet_leaf_121_clk _01295_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11993_ sha256cu.msg_scheduler.mreg_14\[27\] _05808_ VGND VGND VPWR VPWR _05809_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13732_ clknet_leaf_83_clk _00278_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10944_ _04704_ _04809_ _04810_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__o21a_2
X_13663_ clknet_leaf_84_clk _00209_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10875_ _01987_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__clkbuf_4
X_13594_ clknet_leaf_67_clk _00140_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_12614_ _06284_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12545_ _06246_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12476_ sha256cu.m_pad_pars.block_512\[7\]\[4\] _06205_ VGND VGND VPWR VPWR _06210_
+ sky130_fd_sc_hd__and2_1
XANTENNA_5 _01494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14215_ clknet_leaf_28_clk _00761_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11427_ _01920_ _05268_ _05270_ _05150_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__a22o_1
XFILLER_153_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ clknet_leaf_35_clk _00692_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11358_ sha256cu.m_pad_pars.block_512\[61\]\[4\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[4\]
+ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a22o_1
XFILLER_152_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10309_ sha256cu.msg_scheduler.mreg_5\[7\] _04407_ _04412_ _04410_ VGND VGND VPWR
+ VPWR _00627_ sky130_fd_sc_hd__o211a_1
XFILLER_98_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14077_ clknet_leaf_36_clk _00623_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ _04747_ _05130_ _05139_ _01985_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__o211a_2
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13028_ _06504_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__clkbuf_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07520_ _02146_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__inv_2
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07451_ sha256cu.iter_processing.w\[2\] _02078_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07382_ _01913_ _02013_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__or2_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09121_ _03603_ _03605_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__or2_1
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_123_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_148_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09052_ _03538_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__nand2_1
X_08003_ sha256cu.K\[16\] _02615_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__nand2_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09954_ sha256cu.msg_scheduler.mreg_1\[15\] _04202_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__or2_1
X_08905_ _03396_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nand2_1
X_09885_ sha256cu.msg_scheduler.mreg_12\[26\] _04167_ _04168_ _04157_ VGND VGND VPWR
+ VPWR _00441_ sky130_fd_sc_hd__o211a_1
XFILLER_58_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ sha256cu.K\[5\] _03298_ _03297_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__a21o_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ sha256cu.m_out_digest.h_in\[4\] sha256cu.m_out_digest.d_in\[4\] VGND VGND
+ VPWR VPWR _03265_ sky130_fd_sc_hd__or2_1
XANTENNA_406 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _02336_ _02337_ _02338_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__and3_1
X_08698_ _03198_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__nand2_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07649_ sha256cu.m_out_digest.a_in\[29\] VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__buf_4
XFILLER_53_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10660_ sha256cu.msg_scheduler.mreg_10\[30\] _04601_ VGND VGND VPWR VPWR _04613_
+ sky130_fd_sc_hd__or2_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09319_ _03794_ _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10591_ sha256cu.msg_scheduler.mreg_9\[0\] _04567_ _04573_ _04570_ VGND VGND VPWR
+ VPWR _00748_ sky130_fd_sc_hd__o211a_1
XFILLER_22_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_114_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ _03288_ _01949_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__and2_1
X_12261_ _06064_ _06065_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__and2_1
X_14000_ clknet_leaf_56_clk _00546_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11212_ sha256cu.m_pad_pars.block_512\[10\]\[5\] _04963_ _05061_ _05065_ VGND VGND
+ VPWR VPWR _05066_ sky130_fd_sc_hd__a211o_1
XFILLER_134_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12192_ _05998_ _05999_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__nand2_1
X_11143_ sha256cu.m_pad_pars.block_512\[2\]\[0\] _04999_ _05001_ sha256cu.m_pad_pars.block_512\[42\]\[0\]
+ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__a22o_1
Xinput120 hash[207] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_4
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11074_ _04760_ _04775_ sha256cu.m_pad_pars.block_512\[3\]\[7\] VGND VGND VPWR VPWR
+ _04934_ sky130_fd_sc_hd__a21oi_1
Xinput142 hash[227] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_2
X_10025_ sha256cu.msg_scheduler.mreg_1\[13\] _04247_ _04249_ _04250_ VGND VGND VPWR
+ VPWR _00505_ sky130_fd_sc_hd__o211a_1
Xinput131 hash[217] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_4
Xinput153 hash[237] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14902_ clknet_leaf_123_clk _01416_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput164 hash[247] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
Xinput186 hash[36] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput175 hash[26] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput197 hash[46] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14833_ clknet_leaf_2_clk _01347_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11976_ _05790_ _05791_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__nand2_1
XFILLER_91_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14764_ clknet_leaf_8_clk _01278_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13715_ clknet_leaf_61_clk _00261_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14695_ clknet_leaf_8_clk _01209_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10927_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__buf_2
X_13646_ clknet_leaf_74_clk _00192_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10858_ sha256cu.m_pad_pars.add_out3\[3\] _04728_ _04730_ _01971_ _01974_ VGND VGND
+ VPWR VPWR _00858_ sky130_fd_sc_hd__o221a_1
XFILLER_118_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10789_ sha256cu.msg_scheduler.mreg_12\[22\] _04679_ VGND VGND VPWR VPWR _04686_
+ sky130_fd_sc_hd__or2_1
X_13577_ clknet_leaf_81_clk _00123_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_105_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_9_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12528_ _06237_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12459_ sha256cu.m_pad_pars.block_512\[6\]\[4\] _06196_ VGND VGND VPWR VPWR _06201_
+ sky130_fd_sc_hd__and2_1
XFILLER_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14129_ clknet_leaf_34_clk _00675_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06951_ _01601_ _01640_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__or2_1
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09670_ _04043_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__clkbuf_4
X_08621_ sha256cu.m_out_digest.c_in\[5\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[5\]
+ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__o22a_1
XFILLER_94_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06882_ sha256cu.msg_scheduler.counter_iteration\[0\] _01574_ _01575_ sha256cu.iter_processing.rst
+ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__o211a_1
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08552_ _03149_ _03150_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__xnor2_1
X_07503_ sha256cu.m_out_digest.a_in\[25\] _02129_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__xnor2_1
X_08483_ _03043_ _03045_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__or2b_1
X_07434_ sha256cu.K\[1\] _02062_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07365_ _01976_ _01998_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__and2_1
XFILLER_136_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09104_ _03588_ _03589_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__nor2_1
X_07296_ sha256cu.m_pad_pars.add_512_block\[3\] sha256cu.m_pad_pars.add_512_block\[2\]
+ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__or2_2
X_09035_ _03522_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09937_ sha256cu.msg_scheduler.mreg_0\[7\] _04195_ _04200_ _04198_ VGND VGND VPWR
+ VPWR _00467_ sky130_fd_sc_hd__o211a_1
XFILLER_104_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09868_ sha256cu.msg_scheduler.mreg_12\[19\] _04153_ _04158_ _04157_ VGND VGND VPWR
+ VPWR _00434_ sky130_fd_sc_hd__o211a_1
XFILLER_58_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _03263_ _03285_ _03309_ _03314_ _03307_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__a311oi_4
X_09799_ sha256cu.msg_scheduler.mreg_14\[22\] _04106_ VGND VGND VPWR VPWR _04119_
+ sky130_fd_sc_hd__or2_1
XFILLER_18_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_214 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ sha256cu.msg_scheduler.mreg_14\[29\] _05652_ VGND VGND VPWR VPWR _05653_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_203 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _05562_ _05563_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__nor2_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_258 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_236 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10712_ sha256cu.msg_scheduler.mreg_10\[20\] _04633_ _04642_ _04636_ VGND VGND VPWR
+ VPWR _00800_ sky130_fd_sc_hd__o211a_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13500_ sha256cu.K\[26\] _06713_ _06718_ _00054_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__a22o_1
X_11692_ _05492_ _05507_ _05520_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a21o_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ clknet_leaf_9_clk _00994_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10643_ sha256cu.msg_scheduler.mreg_9\[22\] _04594_ _04603_ _04597_ VGND VGND VPWR
+ VPWR _00770_ sky130_fd_sc_hd__o211a_1
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13431_ _03288_ _06720_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__and2_1
X_10574_ sha256cu.msg_scheduler.mreg_9\[25\] _04561_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__or2_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13362_ _06681_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_1
X_12313_ sha256cu.data_in_padd\[30\] _05433_ _05445_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13293_ sha256cu.m_pad_pars.block_512\[55\]\[1\] _06644_ VGND VGND VPWR VPWR _06646_
+ sky130_fd_sc_hd__and2_1
X_12244_ _06024_ _06030_ _06048_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__or3_1
X_12175_ _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__inv_2
X_11126_ sha256cu.m_pad_pars.block_512\[58\]\[0\] _01920_ _04982_ _04983_ _04984_
+ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__a32o_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11057_ _04913_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__buf_4
XFILLER_49_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10008_ sha256cu.msg_scheduler.mreg_1\[6\] _04234_ _04240_ _04237_ VGND VGND VPWR
+ VPWR _00498_ sky130_fd_sc_hd__o211a_1
X_14816_ clknet_leaf_96_clk _01330_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11959_ sha256cu.msg_scheduler.mreg_9\[16\] sha256cu.msg_scheduler.mreg_0\[16\] VGND
+ VGND VPWR VPWR _05776_ sky130_fd_sc_hd__or2_1
X_14747_ clknet_leaf_125_clk _01261_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14678_ clknet_leaf_114_clk _01192_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13629_ clknet_leaf_68_clk _00175_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07150_ _01650_ _01728_ _01819_ _01821_ _01629_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__o311a_1
X_07081_ _00457_ _01755_ _01756_ _01760_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__a31o_1
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07983_ sha256cu.iter_processing.w\[16\] _02596_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__xnor2_1
X_09722_ sha256cu.iter_processing.w\[21\] _04067_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__or2_1
XFILLER_95_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06934_ _01573_ _01577_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__or2_2
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09653_ sha256cu.m_out_digest.h_in\[17\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[17\]
+ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__a22o_1
X_06865_ state\[0\] VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__inv_2
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09584_ sha256cu.m_out_digest.f_in\[24\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[24\]
+ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o22a_1
X_08604_ sha256cu.m_out_digest.b_in\[22\] _03177_ _03176_ _02026_ VGND VGND VPWR VPWR
+ _00149_ sky130_fd_sc_hd__o22a_1
X_06796_ net217 net220 net219 net222 VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__or4_2
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08535_ _03088_ _03089_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__and2b_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08466_ _03035_ _03036_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__o21bai_2
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07417_ _02043_ _02044_ _02045_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__and3_1
X_08397_ sha256cu.m_out_digest.e_in\[6\] sha256cu.m_out_digest.e_in\[1\] VGND VGND
+ VPWR VPWR _03000_ sky130_fd_sc_hd__xnor2_4
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07348_ sha256cu.m_pad_pars.add_out1\[5\] _01984_ _01981_ _01988_ VGND VGND VPWR
+ VPWR _00084_ sky130_fd_sc_hd__a31o_1
XFILLER_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07279_ sha256cu.m_pad_pars.m_size\[3\] sha256cu.m_pad_pars.block_512\[63\]\[3\]
+ _01928_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__mux2_1
XFILLER_152_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10290_ sha256cu.msg_scheduler.mreg_5\[31\] _04401_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__or2_1
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09018_ sha256cu.m_out_digest.h_in\[13\] sha256cu.m_out_digest.d_in\[13\] VGND VGND
+ VPWR VPWR _03507_ sky130_fd_sc_hd__nor2_1
XFILLER_105_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13980_ clknet_leaf_55_clk _00526_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12931_ _06270_ _04995_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__nand2_2
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12862_ _02111_ _05081_ _04975_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__or3_2
XFILLER_46_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _05620_ _05616_ _05634_ _05635_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__nand4_1
XFILLER_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14601_ clknet_leaf_14_clk _01115_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _06379_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__clkbuf_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ sha256cu.msg_scheduler.mreg_9\[7\] sha256cu.msg_scheduler.mreg_0\[7\] VGND
+ VGND VPWR VPWR _05570_ sky130_fd_sc_hd__or2_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ clknet_leaf_106_clk _01046_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11675_ _05502_ _05503_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__a21o_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ clknet_leaf_98_clk _00977_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10626_ sha256cu.msg_scheduler.mreg_9\[15\] _04581_ _04593_ _04584_ VGND VGND VPWR
+ VPWR _00763_ sky130_fd_sc_hd__o211a_1
X_13414_ _06708_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14394_ clknet_leaf_47_clk _00908_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_143_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10557_ _04447_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__buf_2
X_13345_ sha256cu.m_pad_pars.block_512\[58\]\[2\] _06671_ VGND VGND VPWR VPWR _06673_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10488_ sha256cu.msg_scheduler.mreg_7\[20\] _04513_ _04514_ _04503_ VGND VGND VPWR
+ VPWR _00704_ sky130_fd_sc_hd__o211a_1
X_13276_ sha256cu.m_pad_pars.block_512\[54\]\[1\] _06635_ VGND VGND VPWR VPWR _06637_
+ sky130_fd_sc_hd__and2_1
X_12227_ sha256cu.msg_scheduler.mreg_9\[27\] sha256cu.msg_scheduler.mreg_0\[27\] VGND
+ VGND VPWR VPWR _06033_ sky130_fd_sc_hd__or2_1
XFILLER_151_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12158_ _05963_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__and2_1
XFILLER_2_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12089_ _05867_ _05871_ _05868_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__a21boi_1
XFILLER_68_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11109_ _04951_ _04967_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__nand2_1
XFILLER_49_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08320_ _02899_ _02896_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__or2b_1
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08251_ sha256cu.m_out_digest.b_in\[23\] sha256cu.m_out_digest.a_in\[23\] _02857_
+ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07202_ _01600_ _01682_ _01694_ _01649_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__a211o_1
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08182_ _02788_ _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07133_ _01632_ _01584_ _01673_ _01805_ _01806_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__o311a_1
XFILLER_146_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07064_ _01626_ _01744_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__nor2_1
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07966_ _02578_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__xor2_2
X_09705_ sha256cu.msg_scheduler.mreg_14\[13\] _04060_ _04065_ _04064_ VGND VGND VPWR
+ VPWR _00364_ sky130_fd_sc_hd__o211a_1
XFILLER_56_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06917_ _01607_ _01608_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__nor2_2
X_07897_ _02481_ _02479_ _02513_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__o21ai_1
X_09636_ _02515_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__buf_4
XFILLER_56_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06848_ net252 net255 net254 net3 VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__or4_1
X_09567_ sha256cu.m_out_digest.f_in\[9\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[9\]
+ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__a22o_1
X_06779_ net34 net67 net56 net89 VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__or4_1
XFILLER_82_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08518_ sha256cu.m_out_digest.e_in\[9\] sha256cu.m_out_digest.e_in\[4\] VGND VGND
+ VPWR VPWR _03118_ sky130_fd_sc_hd__xnor2_4
X_09498_ _03965_ _03969_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__and2_1
XFILLER_70_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08449_ sha256cu.m_out_digest.b_in\[28\] _02232_ _03050_ VGND VGND VPWR VPWR _03051_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11460_ _04760_ _04801_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__a21oi_1
X_10411_ sha256cu.msg_scheduler.mreg_7\[19\] _04468_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__or2_1
XFILLER_99_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11391_ _01952_ _05233_ _05234_ sha256cu.m_pad_pars.block_512\[53\]\[7\] VGND VGND
+ VPWR VPWR _05235_ sky130_fd_sc_hd__o22a_1
XFILLER_152_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10342_ sha256cu.msg_scheduler.mreg_5\[21\] _04421_ _04431_ _04424_ VGND VGND VPWR
+ VPWR _00641_ sky130_fd_sc_hd__o211a_1
X_13130_ sha256cu.m_pad_pars.block_512\[45\]\[5\] _06553_ VGND VGND VPWR VPWR _06559_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13061_ sha256cu.m_pad_pars.block_512\[41\]\[5\] _06516_ VGND VGND VPWR VPWR _06522_
+ sky130_fd_sc_hd__and2_1
X_10273_ sha256cu.msg_scheduler.mreg_4\[24\] _04380_ _04391_ _04383_ VGND VGND VPWR
+ VPWR _00612_ sky130_fd_sc_hd__o211a_1
X_12012_ _05798_ _05802_ _05799_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a21boi_1
XFILLER_105_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13963_ clknet_leaf_55_clk _00509_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_74_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_85_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13894_ clknet_leaf_24_clk _00440_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12914_ _01912_ _05146_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__or2_2
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12845_ _06251_ _05081_ _05124_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__or3_4
XFILLER_34_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12776_ _06370_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__clkbuf_1
X_11727_ sha256cu.msg_scheduler.mreg_1\[24\] _05553_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__xnor2_2
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ clknet_leaf_4_clk _01029_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11658_ sha256cu.msg_scheduler.mreg_1\[10\] sha256cu.msg_scheduler.mreg_1\[6\] VGND
+ VGND VPWR VPWR _05488_ sky130_fd_sc_hd__xnor2_1
X_14446_ clknet_leaf_112_clk _00960_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10609_ sha256cu.msg_scheduler.mreg_9\[7\] _04581_ _04583_ _04584_ VGND VGND VPWR
+ VPWR _00755_ sky130_fd_sc_hd__o211a_1
X_14377_ clknet_leaf_110_clk _00891_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11589_ _05315_ _05424_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__or2b_1
XFILLER_116_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13328_ sha256cu.m_pad_pars.block_512\[57\]\[2\] _06660_ VGND VGND VPWR VPWR _06664_
+ sky130_fd_sc_hd__and2_1
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13259_ sha256cu.m_pad_pars.block_512\[53\]\[1\] _06626_ VGND VGND VPWR VPWR _06628_
+ sky130_fd_sc_hd__and2_1
XFILLER_124_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07820_ _02064_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__clkbuf_4
X_07751_ sha256cu.iter_processing.w\[9\] _02340_ _02339_ VGND VGND VPWR VPWR _02371_
+ sky130_fd_sc_hd__a21o_1
XFILLER_84_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_76_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_38_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07682_ sha256cu.m_out_digest.a_in\[30\] VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__buf_4
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09421_ _03839_ _03895_ _03896_ _03893_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__o211ai_1
XFILLER_64_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09352_ _03828_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__xor2_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08303_ _02907_ _02908_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__or2_1
XFILLER_138_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09283_ _03760_ _03761_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__and2_1
XFILLER_33_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08234_ _02798_ _02800_ _02841_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08165_ sha256cu.m_out_digest.a_in\[23\] _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07116_ _01637_ _01642_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__nand2_1
XFILLER_134_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08096_ sha256cu.m_out_digest.b_in\[19\] _02233_ _02706_ VGND VGND VPWR VPWR _02707_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07047_ _01609_ _01726_ _01728_ _01655_ _01729_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__o32a_1
XFILLER_133_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08998_ _03486_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__nor2_1
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_67_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
X_07949_ sha256cu.m_out_digest.e_in\[21\] sha256cu.m_out_digest.e_in\[8\] VGND VGND
+ VPWR VPWR _02564_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10960_ _04705_ _04770_ _04807_ _04746_ _04771_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__o32a_1
X_09619_ _02112_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__buf_4
X_10891_ _01940_ _04752_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__or2_2
XFILLER_71_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12630_ sha256cu.m_pad_pars.block_512\[16\]\[3\] _06289_ VGND VGND VPWR VPWR _06293_
+ sky130_fd_sc_hd__and2_1
X_12561_ sha256cu.m_pad_pars.block_512\[12\]\[3\] _06252_ VGND VGND VPWR VPWR _06256_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12492_ _06218_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__clkbuf_1
X_14300_ clknet_leaf_95_clk _00022_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__dfxtp_1
X_11512_ sha256cu.m_pad_pars.block_512\[28\]\[3\] _05296_ _05351_ _01921_ VGND VGND
+ VPWR VPWR _05352_ sky130_fd_sc_hd__a22o_1
XFILLER_109_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14231_ clknet_leaf_27_clk _00777_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11443_ _04808_ _04819_ _04824_ _05264_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__o22a_1
X_14162_ clknet_leaf_34_clk _00708_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11374_ _05212_ _05214_ _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__or3_1
X_13113_ sha256cu.m_pad_pars.block_512\[44\]\[5\] _06544_ VGND VGND VPWR VPWR _06550_
+ sky130_fd_sc_hd__and2_1
X_14093_ clknet_leaf_32_clk _00639_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10325_ sha256cu.msg_scheduler.mreg_6\[14\] _04415_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__or2_1
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10256_ sha256cu.msg_scheduler.mreg_5\[17\] _04374_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__or2_1
XFILLER_79_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13044_ sha256cu.m_pad_pars.block_512\[40\]\[5\] _06507_ VGND VGND VPWR VPWR _06513_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10187_ sha256cu.msg_scheduler.mreg_4\[19\] _04335_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__or2_1
XFILLER_94_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_58_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_47_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_13946_ clknet_leaf_43_clk _00492_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13877_ clknet_leaf_20_clk _00423_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12828_ _06251_ _05081_ _05295_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__or3_2
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _06361_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14429_ clknet_leaf_119_clk _00943_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09970_ sha256cu.msg_scheduler.mreg_1\[22\] _04215_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__or2_1
XFILLER_89_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08921_ _03394_ _03395_ _03412_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__and3_1
XFILLER_131_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08852_ _03345_ _03346_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__nand2_1
X_07803_ _02418_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__xnor2_2
XFILLER_112_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08783_ _03264_ _03279_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_49_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_85_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07734_ _02300_ _02311_ _02354_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__o21ba_1
X_07665_ _02285_ _02287_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__xor2_2
XFILLER_38_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09404_ _03878_ _03879_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__nor2_1
XFILLER_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07596_ _02037_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ sha256cu.m_out_digest.h_in\[24\] sha256cu.m_out_digest.d_in\[24\] VGND VGND
+ VPWR VPWR _03813_ sky130_fd_sc_hd__or2_1
XFILLER_139_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09266_ sha256cu.K\[20\] _03706_ _03705_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__a21o_1
X_08217_ _02778_ _02781_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__nand2_1
X_09197_ sha256cu.K\[19\] _03679_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__xor2_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08148_ sha256cu.K\[20\] _02757_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__xnor2_2
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08079_ _02666_ _02690_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__xnor2_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10110_ sha256cu.msg_scheduler.mreg_3\[18\] _04295_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__or2_1
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11090_ _04736_ _04764_ _04932_ _04941_ _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__a311o_1
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10041_ sha256cu.msg_scheduler.mreg_2\[21\] _04254_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__or2_1
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11992_ sha256cu.msg_scheduler.mreg_14\[4\] sha256cu.msg_scheduler.mreg_14\[2\] VGND
+ VGND VPWR VPWR _05808_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13800_ clknet_leaf_81_clk _00346_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14780_ clknet_leaf_126_clk _01294_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13731_ clknet_leaf_83_clk _00277_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10943_ sha256cu.m_pad_pars.add_out3\[3\] sha256cu.m_pad_pars.add_out3\[2\] _04756_
+ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__and3_1
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13662_ clknet_leaf_69_clk _00208_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10874_ _01980_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13593_ clknet_leaf_64_clk _00139_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12613_ sha256cu.m_pad_pars.block_512\[15\]\[3\] _06280_ VGND VGND VPWR VPWR _06284_
+ sky130_fd_sc_hd__and2_1
XFILLER_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12544_ sha256cu.m_pad_pars.block_512\[11\]\[4\] _06241_ VGND VGND VPWR VPWR _06246_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12475_ _06209_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14214_ clknet_leaf_27_clk _00760_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_6 _01494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11426_ _01950_ _05136_ _05269_ sha256cu.m_pad_pars.block_512\[49\]\[7\] VGND VGND
+ VPWR VPWR _05270_ sky130_fd_sc_hd__o22a_1
X_14145_ clknet_leaf_35_clk _00691_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11357_ sha256cu.m_pad_pars.block_512\[1\]\[4\] _05135_ _05158_ sha256cu.m_pad_pars.block_512\[21\]\[4\]
+ _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__a221o_1
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10308_ sha256cu.msg_scheduler.mreg_6\[7\] _04401_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__or2_1
X_14076_ clknet_leaf_36_clk _00622_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13027_ sha256cu.m_pad_pars.block_512\[39\]\[5\] _06498_ VGND VGND VPWR VPWR _06504_
+ sky130_fd_sc_hd__and2_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ sha256cu.m_pad_pars.add_out1\[2\] sha256cu.m_pad_pars.add_out1\[3\] VGND
+ VGND VPWR VPWR _05139_ sky130_fd_sc_hd__and2b_2
X_10239_ sha256cu.msg_scheduler.mreg_4\[9\] _04367_ _04372_ _04370_ VGND VGND VPWR
+ VPWR _00597_ sky130_fd_sc_hd__o211a_1
XFILLER_79_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13929_ clknet_leaf_52_clk _00475_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_07450_ _02076_ _02077_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__and2b_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07381_ sha256cu.m_out_digest.H7\[0\] _02011_ _02009_ VGND VGND VPWR VPWR _02013_
+ sky130_fd_sc_hd__mux2_1
X_09120_ _03603_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__nand2_1
XFILLER_148_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09051_ _03536_ _03537_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__nand2_1
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08002_ sha256cu.K\[16\] _02615_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__or2_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09953_ sha256cu.msg_scheduler.mreg_0\[14\] _04208_ _04209_ _04198_ VGND VGND VPWR
+ VPWR _00474_ sky130_fd_sc_hd__o211a_1
X_08904_ sha256cu.m_out_digest.h_in\[9\] sha256cu.m_out_digest.d_in\[9\] VGND VGND
+ VPWR VPWR _03397_ sky130_fd_sc_hd__nand2_1
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09884_ sha256cu.msg_scheduler.mreg_13\[26\] _04160_ VGND VGND VPWR VPWR _04168_
+ sky130_fd_sc_hd__or2_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _03329_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__and2_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ sha256cu.K\[3\] _03242_ _03241_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a21bo_1
XFILLER_100_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ sha256cu.m_out_digest.g_in\[9\] sha256cu.m_out_digest.f_in\[9\] sha256cu.m_out_digest.e_in\[9\]
+ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__mux2_1
XANTENNA_407 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ sha256cu.m_out_digest.h_in\[0\] sha256cu.m_out_digest.d_in\[0\] VGND VGND
+ VPWR VPWR _03199_ sky130_fd_sc_hd__or2_1
XFILLER_14_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07648_ _02270_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__inv_2
XFILLER_26_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07579_ _02160_ _02165_ _02203_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__o21a_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09318_ _03795_ _03796_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__nand2_1
XFILLER_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10590_ sha256cu.msg_scheduler.mreg_10\[0\] _04561_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__or2_1
XFILLER_108_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09249_ sha256cu.m_out_digest.h_in\[21\] sha256cu.m_out_digest.d_in\[21\] VGND VGND
+ VPWR VPWR _03730_ sky130_fd_sc_hd__nand2_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12260_ _06062_ _06063_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nand2_1
XFILLER_135_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12191_ sha256cu.msg_scheduler.mreg_14\[12\] sha256cu.msg_scheduler.mreg_14\[10\]
+ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__xor2_1
X_11211_ sha256cu.m_pad_pars.block_512\[6\]\[5\] _04957_ _05001_ sha256cu.m_pad_pars.block_512\[42\]\[5\]
+ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__a221o_1
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11142_ _04721_ _04958_ _05000_ _04725_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__and4b_4
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 hash[199] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_2
XFILLER_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11073_ _04769_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__buf_4
X_10024_ _04116_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__buf_2
Xinput154 hash[238] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput132 hash[218] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_4
Xinput143 hash[228] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput121 hash[208] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
X_14901_ clknet_leaf_124_clk _01415_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput187 hash[37] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
Xinput176 hash[27] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput165 hash[248] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14832_ clknet_leaf_4_clk _01346_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput198 hash[47] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
X_11975_ _05790_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__or2_1
X_14763_ clknet_leaf_11_clk _01277_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13714_ clknet_leaf_60_clk _00260_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14694_ clknet_leaf_116_clk _01208_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10926_ _04703_ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__or2_1
X_13645_ clknet_leaf_71_clk _00191_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10857_ sha256cu.m_pad_pars.add_out3\[3\] sha256cu.m_pad_pars.add_out3\[2\] VGND
+ VGND VPWR VPWR _04730_ sky130_fd_sc_hd__nand2_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ _04580_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__clkbuf_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ clknet_leaf_86_clk _00122_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[27\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12527_ sha256cu.m_pad_pars.block_512\[10\]\[4\] _06232_ VGND VGND VPWR VPWR _06237_
+ sky130_fd_sc_hd__and2_1
XFILLER_9_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12458_ _06200_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11409_ _01985_ _05139_ _05243_ _05245_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__a311o_1
X_12389_ sha256cu.m_pad_pars.block_512\[2\]\[3\] _06160_ VGND VGND VPWR VPWR _06164_
+ sky130_fd_sc_hd__and2_1
X_14128_ clknet_leaf_33_clk _00674_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14059_ clknet_leaf_39_clk _00605_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06950_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__clkbuf_4
XFILLER_140_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06881_ sha256cu.counter_iteration\[0\] _01568_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__or2_1
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08620_ sha256cu.m_out_digest.c_in\[4\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[4\]
+ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__o22a_1
XFILLER_67_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08551_ _03134_ _03136_ _03132_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__o21a_1
X_07502_ _02128_ sha256cu.m_out_digest.a_in\[5\] VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__xnor2_1
X_08482_ _03080_ _03082_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__xnor2_1
X_07433_ _02042_ _02061_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09103_ _02565_ _03561_ _03562_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__a21boi_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07364_ sha256cu.m_pad_pars.add_out0\[5\] _01993_ _01999_ _02000_ VGND VGND VPWR
+ VPWR _00088_ sky130_fd_sc_hd__o211a_1
XFILLER_149_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07295_ sha256cu.m_pad_pars.add_512_block\[0\] VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__clkbuf_4
X_09034_ sha256cu.K\[12\] _03484_ _03483_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a21o_1
XFILLER_132_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09936_ sha256cu.msg_scheduler.mreg_1\[7\] _04174_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__or2_1
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09867_ sha256cu.msg_scheduler.mreg_13\[19\] _04147_ VGND VGND VPWR VPWR _04158_
+ sky130_fd_sc_hd__or2_1
XFILLER_19_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _03282_ _03284_ _03308_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__nor3_1
XFILLER_93_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09798_ sha256cu.msg_scheduler.mreg_13\[21\] _04112_ _04118_ _04117_ VGND VGND VPWR
+ VPWR _00404_ sky130_fd_sc_hd__o211a_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_215 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _02126_ _03247_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__xor2_1
XFILLER_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_204 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _05562_ _05563_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__nand2_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_248 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_237 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_226 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10711_ sha256cu.msg_scheduler.mreg_11\[20\] _04640_ VGND VGND VPWR VPWR _04642_
+ sky130_fd_sc_hd__or2_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11691_ _05517_ _05519_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__xnor2_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10642_ sha256cu.msg_scheduler.mreg_10\[22\] _04601_ VGND VGND VPWR VPWR _04603_
+ sky130_fd_sc_hd__or2_1
XFILLER_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13430_ sha256cu.K\[0\] _06714_ _06719_ _00036_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__a22o_1
XFILLER_139_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10573_ sha256cu.msg_scheduler.mreg_8\[24\] _04554_ _04563_ _04557_ VGND VGND VPWR
+ VPWR _00740_ sky130_fd_sc_hd__o211a_1
XFILLER_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13361_ sha256cu.m_pad_pars.block_512\[59\]\[2\] _06671_ VGND VGND VPWR VPWR _06681_
+ sky130_fd_sc_hd__and2_1
X_12312_ _06112_ _06114_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__nand2_1
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13292_ _06645_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
X_12243_ _06024_ _06030_ _06048_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12174_ _05981_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__and2_1
XFILLER_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11125_ sha256cu.m_pad_pars.add_out2\[5\] sha256cu.m_pad_pars.add_out2\[4\] sha256cu.m_pad_pars.add_out2\[3\]
+ sha256cu.m_pad_pars.add_out2\[2\] VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__and4_2
XFILLER_110_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11056_ _04810_ _04911_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__a21o_1
X_10007_ sha256cu.msg_scheduler.mreg_2\[6\] _04228_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__or2_1
XFILLER_49_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14815_ clknet_leaf_98_clk _01329_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14746_ clknet_leaf_125_clk _01260_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11958_ _05747_ _05750_ _05769_ _05768_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__a31oi_4
XFILLER_60_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11889_ sha256cu.data_in_padd\[12\] _05433_ _05707_ _05709_ _04046_ VGND VGND VPWR
+ VPWR _05710_ sky130_fd_sc_hd__a221o_1
X_10909_ sha256cu.m_pad_pars.add_512_block\[3\] sha256cu.m_pad_pars.add_512_block\[2\]
+ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__nand2_2
XFILLER_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14677_ clknet_leaf_1_clk _01191_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13628_ clknet_leaf_68_clk _00174_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13559_ clknet_leaf_63_clk _00105_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_146_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07080_ _01758_ _01759_ _01631_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a21oi_1
XFILLER_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07982_ _02594_ _02595_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09721_ sha256cu.msg_scheduler.mreg_14\[20\] _04073_ _04074_ _04064_ VGND VGND VPWR
+ VPWR _00371_ sky130_fd_sc_hd__o211a_1
X_06933_ _01622_ _01623_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__nor2_1
XFILLER_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09652_ sha256cu.m_out_digest.h_in\[16\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[16\]
+ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__a22o_1
X_06864_ net257 _01561_ state\[1\] VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__nor3b_1
XFILLER_94_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09583_ sha256cu.m_out_digest.f_in\[23\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[23\]
+ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__a22o_1
X_06795_ net208 net211 net210 net214 VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__or4_2
X_08603_ sha256cu.m_out_digest.b_in\[21\] _03177_ _03176_ sha256cu.m_out_digest.a_in\[21\]
+ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__o22a_1
XFILLER_83_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08534_ _03132_ _03133_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__nand2_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08465_ _03037_ _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07416_ sha256cu.m_out_digest.g_in\[1\] sha256cu.m_out_digest.f_in\[1\] sha256cu.m_out_digest.e_in\[1\]
+ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__mux2_1
X_08396_ sha256cu.m_out_digest.h_in\[27\] _02998_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07347_ _01977_ _01985_ _01987_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__and3_1
XFILLER_149_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09017_ _03479_ _03480_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nor2_1
X_07278_ _01923_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09919_ sha256cu.msg_scheduler.temp_case _04190_ _02000_ VGND VGND VPWR VPWR _00459_
+ sky130_fd_sc_hd__o21a_1
XFILLER_92_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12930_ _06452_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__clkbuf_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _06415_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__clkbuf_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _05620_ _05616_ _05634_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__a22o_1
XFILLER_73_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14600_ clknet_leaf_14_clk _01114_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12792_ sha256cu.m_pad_pars.block_512\[25\]\[7\] _05243_ _06351_ VGND VGND VPWR VPWR
+ _06379_ sky130_fd_sc_hd__mux2_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ sha256cu.iter_processing.w\[6\] _05430_ _05569_ _05335_ VGND VGND VPWR VPWR
+ _00904_ sky130_fd_sc_hd__o211a_1
X_14531_ clknet_leaf_106_clk _01045_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ sha256cu.data_in_padd\[3\] _05447_ _04692_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__a21o_1
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14462_ clknet_leaf_115_clk _00976_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10625_ sha256cu.msg_scheduler.mreg_10\[15\] _04588_ VGND VGND VPWR VPWR _04593_
+ sky130_fd_sc_hd__or2_1
X_13413_ sha256cu.m_pad_pars.block_512\[62\]\[3\] _01928_ VGND VGND VPWR VPWR _06708_
+ sky130_fd_sc_hd__and2_1
XFILLER_128_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14393_ clknet_leaf_47_clk _00907_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10556_ sha256cu.msg_scheduler.mreg_8\[17\] _04540_ _04553_ _04543_ VGND VGND VPWR
+ VPWR _00733_ sky130_fd_sc_hd__o211a_1
X_13344_ _06672_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10487_ sha256cu.msg_scheduler.mreg_8\[20\] _04507_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__or2_1
X_13275_ _06636_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12226_ sha256cu.iter_processing.w\[26\] _05894_ _06032_ _05866_ VGND VGND VPWR VPWR
+ _00924_ sky130_fd_sc_hd__o211a_1
X_12157_ _05889_ _05961_ _05964_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__o211a_1
XFILLER_69_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11108_ _04966_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__inv_2
XFILLER_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12088_ _05897_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__xor2_1
XFILLER_96_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11039_ sha256cu.m_pad_pars.block_512\[39\]\[6\] _04800_ _04831_ sha256cu.m_pad_pars.block_512\[19\]\[6\]
+ _04899_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__a221o_1
XFILLER_49_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14729_ clknet_leaf_7_clk _01243_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08250_ sha256cu.m_out_digest.b_in\[23\] sha256cu.m_out_digest.a_in\[23\] sha256cu.m_out_digest.c_in\[23\]
+ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__a21o_1
XFILLER_33_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08181_ _02742_ _02751_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a21oi_1
X_07201_ _00455_ _01696_ _01689_ _01585_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__a211o_1
X_07132_ _01667_ _01583_ _01640_ _01570_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__o31a_1
XFILLER_146_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07063_ _01743_ _01646_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__nand2_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07965_ _02518_ _02537_ _02579_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__a21oi_2
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09704_ sha256cu.iter_processing.w\[13\] _04054_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__or2_1
X_06916_ _01577_ _01600_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__nor2_8
X_07896_ _02511_ _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nor2_1
X_09635_ sha256cu.m_out_digest.h_in\[2\] _04037_ _04036_ sha256cu.m_out_digest.g_in\[2\]
+ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__a22o_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06847_ net243 net247 net246 net249 VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__or4_2
X_09566_ sha256cu.m_out_digest.f_in\[8\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[8\]
+ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__a22o_1
XFILLER_82_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06778_ net112 net190 net179 net212 VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__or4_2
X_08517_ sha256cu.m_out_digest.h_in\[30\] _03116_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__xnor2_1
X_09497_ _03965_ _03969_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__nor2_1
XFILLER_142_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08448_ sha256cu.m_out_digest.b_in\[28\] _02232_ sha256cu.m_out_digest.c_in\[28\]
+ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__a21o_1
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10410_ sha256cu.msg_scheduler.mreg_6\[18\] _04461_ _04470_ _04464_ VGND VGND VPWR
+ VPWR _00670_ sky130_fd_sc_hd__o211a_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08379_ _02981_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__or2b_1
XFILLER_11_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ _04824_ _04969_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__nor2_1
XFILLER_152_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10341_ sha256cu.msg_scheduler.mreg_6\[21\] _04428_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__or2_1
XFILLER_137_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10272_ sha256cu.msg_scheduler.mreg_5\[24\] _04387_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__or2_1
X_13060_ _06521_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12011_ _05823_ _05825_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__xor2_1
XFILLER_79_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13962_ clknet_leaf_59_clk _00508_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12913_ _06443_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__clkbuf_1
X_13893_ clknet_leaf_24_clk _00439_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12844_ _06406_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__clkbuf_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ sha256cu.m_pad_pars.block_512\[24\]\[7\] _05405_ _06351_ VGND VGND VPWR VPWR
+ _06370_ sky130_fd_sc_hd__mux2_1
X_11726_ sha256cu.msg_scheduler.mreg_1\[13\] sha256cu.msg_scheduler.mreg_1\[9\] VGND
+ VGND VPWR VPWR _05553_ sky130_fd_sc_hd__xnor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14514_ clknet_leaf_4_clk _01028_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11657_ _05485_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__nand2_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14445_ clknet_leaf_8_clk _00959_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10608_ _04529_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__buf_2
X_14376_ clknet_leaf_110_clk _00890_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_11588_ _04786_ _04924_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10539_ sha256cu.msg_scheduler.mreg_9\[10\] _04534_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__or2_1
X_13327_ _06663_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13258_ _06627_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
X_12209_ _05989_ _05993_ _05990_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__a21boi_1
XFILLER_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13189_ sha256cu.m_pad_pars.block_512\[49\]\[0\] _06590_ VGND VGND VPWR VPWR _06591_
+ sky130_fd_sc_hd__and2_1
X_07750_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__buf_4
XFILLER_84_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07681_ _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__inv_2
XFILLER_92_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09420_ _03863_ _03869_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__or2_1
XFILLER_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09351_ _03794_ _03797_ _03796_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09282_ _03760_ _03761_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__nor2_1
X_08302_ _02889_ _02890_ _02906_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__and3_1
XFILLER_21_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08233_ _02798_ _02800_ _02758_ _02760_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a211o_1
XFILLER_20_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08164_ sha256cu.m_out_digest.a_in\[11\] sha256cu.m_out_digest.a_in\[2\] VGND VGND
+ VPWR VPWR _02773_ sky130_fd_sc_hd__xnor2_2
XFILLER_134_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08095_ sha256cu.m_out_digest.b_in\[19\] _02233_ sha256cu.m_out_digest.c_in\[19\]
+ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__a21o_1
X_07115_ _01578_ _01690_ _01703_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__a31o_1
X_07046_ _01607_ _01606_ _01588_ _01583_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__a31o_1
XFILLER_134_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08997_ _03481_ _03485_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__and2_1
X_07948_ sha256cu.iter_processing.w\[15\] _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__xnor2_2
X_07879_ sha256cu.m_out_digest.h_in\[13\] _02495_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09618_ sha256cu.m_out_digest.g_in\[20\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[20\]
+ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__a22o_1
XFILLER_55_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10890_ _04747_ _04754_ _04755_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__o211a_2
X_09549_ _04018_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ _06255_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__clkbuf_1
X_12491_ sha256cu.m_pad_pars.block_512\[8\]\[3\] _06214_ VGND VGND VPWR VPWR _06218_
+ sky130_fd_sc_hd__and2_1
X_11511_ sha256cu.m_pad_pars.block_512\[60\]\[3\] _01998_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[3\]
+ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__a22o_1
XFILLER_109_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14230_ clknet_leaf_27_clk _00776_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11442_ _01935_ _05277_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__and3_2
XFILLER_153_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14161_ clknet_leaf_34_clk _00707_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11373_ sha256cu.m_pad_pars.block_512\[9\]\[5\] _05144_ _05147_ sha256cu.m_pad_pars.block_512\[33\]\[5\]
+ _05218_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__a221o_1
X_10324_ _04314_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__buf_2
X_13112_ _06549_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__clkbuf_1
X_14092_ clknet_leaf_37_clk _00638_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10255_ sha256cu.msg_scheduler.mreg_4\[16\] _04380_ _04381_ _04370_ VGND VGND VPWR
+ VPWR _00604_ sky130_fd_sc_hd__o211a_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _06512_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__clkbuf_1
X_10186_ sha256cu.msg_scheduler.mreg_3\[18\] _04341_ _04342_ _04331_ VGND VGND VPWR
+ VPWR _00574_ sky130_fd_sc_hd__o211a_1
XFILLER_121_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13945_ clknet_leaf_43_clk _00491_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13876_ clknet_leaf_20_clk _00422_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12827_ _06397_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ sha256cu.m_pad_pars.block_512\[23\]\[7\] _04927_ _06351_ VGND VGND VPWR VPWR
+ _06361_ sky130_fd_sc_hd__mux2_1
X_11709_ _05535_ _05536_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__nor2_1
X_12689_ sha256cu.m_pad_pars.block_512\[19\]\[7\] _04943_ _06249_ VGND VGND VPWR VPWR
+ _06324_ sky130_fd_sc_hd__mux2_1
X_14428_ clknet_leaf_117_clk _00942_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14359_ clknet_leaf_14_clk _00873_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_08920_ _03394_ _03395_ _03412_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08851_ sha256cu.iter_processing.w\[7\] _02264_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__or2_1
XFILLER_97_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07802_ sha256cu.m_out_digest.h_in\[11\] _02420_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__xnor2_2
X_08782_ _03264_ _03279_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__nand2_1
XFILLER_97_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07733_ _02308_ _02310_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__nor2_1
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07664_ _02221_ _02244_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__a21oi_2
XFILLER_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09403_ sha256cu.iter_processing.w\[26\] _02971_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__and2_1
X_07595_ _02219_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09334_ _03810_ _03811_ _03812_ _03366_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__o211a_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09265_ _03744_ _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__and2_1
X_09196_ _03677_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__nand2_1
X_08216_ _02816_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08147_ _02735_ _02756_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__xnor2_2
XFILLER_106_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08078_ _02688_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__or2_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07029_ _01598_ _01689_ _01711_ _01712_ _01618_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__o32a_1
X_10040_ sha256cu.msg_scheduler.mreg_1\[20\] _04247_ _04258_ _04250_ VGND VGND VPWR
+ VPWR _00512_ sky130_fd_sc_hd__o211a_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11991_ _05805_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__nor2_1
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13730_ clknet_leaf_83_clk _00276_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10942_ _04805_ _04779_ _04807_ _04808_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__o22a_1
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13661_ clknet_leaf_68_clk _00207_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10873_ sha256cu.flag_0_15 _01966_ _01938_ _00896_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__a22o_1
XFILLER_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13592_ clknet_leaf_63_clk _00138_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12612_ _06283_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12543_ _06245_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14213_ clknet_leaf_28_clk _00759_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12474_ sha256cu.m_pad_pars.block_512\[7\]\[3\] _06205_ VGND VGND VPWR VPWR _06209_
+ sky130_fd_sc_hd__and2_1
XANTENNA_7 _01509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11425_ _04824_ _05004_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__nor2_1
XFILLER_153_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14144_ clknet_leaf_35_clk _00690_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11356_ sha256cu.m_pad_pars.block_512\[17\]\[4\] _05138_ _05151_ sha256cu.m_pad_pars.block_512\[49\]\[4\]
+ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__a22o_1
X_10307_ sha256cu.msg_scheduler.mreg_5\[6\] _04407_ _04411_ _04410_ VGND VGND VPWR
+ VPWR _00626_ sky130_fd_sc_hd__o211a_1
X_14075_ clknet_leaf_44_clk _00621_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13026_ _06503_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__clkbuf_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _01985_ _05134_ _05137_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__and3_2
X_10238_ sha256cu.msg_scheduler.mreg_5\[9\] _04361_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__or2_1
X_10169_ sha256cu.msg_scheduler.mreg_4\[11\] _04322_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__or2_1
XFILLER_120_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13928_ clknet_leaf_53_clk _00474_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13859_ clknet_leaf_23_clk _00405_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07380_ sha256cu.m_out_digest.temp_delay _02009_ _02000_ VGND VGND VPWR VPWR _00092_
+ sky130_fd_sc_hd__o21a_1
XFILLER_16_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09050_ _03536_ _03537_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__or2_1
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08001_ _02612_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09952_ sha256cu.msg_scheduler.mreg_1\[14\] _04202_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__or2_1
XFILLER_143_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08903_ sha256cu.m_out_digest.h_in\[9\] sha256cu.m_out_digest.d_in\[9\] VGND VGND
+ VPWR VPWR _03396_ sky130_fd_sc_hd__or2_1
XFILLER_106_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09883_ _04166_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _03316_ _03317_ _03328_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__or3_1
XFILLER_112_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _03237_ _03258_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a21o_1
XFILLER_100_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ sha256cu.m_out_digest.b_in\[9\] sha256cu.m_out_digest.a_in\[9\] sha256cu.m_out_digest.c_in\[9\]
+ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__a21o_1
XFILLER_72_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_408 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ sha256cu.m_out_digest.h_in\[0\] sha256cu.m_out_digest.d_in\[0\] VGND VGND
+ VPWR VPWR _03198_ sky130_fd_sc_hd__nand2_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07647_ sha256cu.m_out_digest.e_in\[18\] _02269_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__xnor2_2
XFILLER_26_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07578_ sha256cu.m_out_digest.h_in\[4\] _02164_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__nand2_1
X_09317_ sha256cu.iter_processing.w\[23\] _02859_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__nand2_1
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09248_ sha256cu.m_out_digest.h_in\[21\] sha256cu.m_out_digest.d_in\[21\] VGND VGND
+ VPWR VPWR _03729_ sky130_fd_sc_hd__or2_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_119_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09179_ _03630_ _03642_ _03661_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__and3_1
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12190_ _05996_ _05997_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__and2_1
X_11210_ sha256cu.m_pad_pars.block_512\[2\]\[5\] _04999_ _04989_ sha256cu.m_pad_pars.block_512\[14\]\[5\]
+ _05063_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__a221o_1
XFILLER_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11141_ _04912_ _04961_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__or2_1
X_11072_ sha256cu.m_pad_pars.block_512\[51\]\[7\] _04825_ _04823_ VGND VGND VPWR VPWR
+ _04932_ sky130_fd_sc_hd__o21ba_1
Xinput100 hash[18] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
Xinput111 hash[19] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput133 hash[219] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_2
X_10023_ sha256cu.msg_scheduler.mreg_2\[13\] _04241_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__or2_1
Xinput144 hash[229] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput122 hash[209] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
X_14900_ clknet_leaf_1_clk _01414_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput166 hash[249] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput177 hash[28] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
Xinput155 hash[239] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_2
X_14831_ clknet_leaf_1_clk _01345_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput199 hash[48] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_4
Xinput188 hash[38] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11974_ _05764_ _05766_ _05762_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__a21oi_1
X_14762_ clknet_leaf_17_clk _01276_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13713_ clknet_leaf_65_clk _00259_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14693_ clknet_leaf_104_clk _01207_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10925_ sha256cu.m_pad_pars.temp_chk _04791_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__or2_2
X_13644_ clknet_leaf_71_clk _00190_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10856_ _04728_ _04729_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__nor2_1
XFILLER_32_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10787_ sha256cu.msg_scheduler.mreg_11\[21\] _04672_ _04684_ _04675_ VGND VGND VPWR
+ VPWR _00833_ sky130_fd_sc_hd__o211a_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ clknet_leaf_86_clk _00121_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12526_ _06236_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12457_ sha256cu.m_pad_pars.block_512\[6\]\[3\] _06196_ VGND VGND VPWR VPWR _06200_
+ sky130_fd_sc_hd__and2_1
X_11408_ _05125_ _05152_ _05247_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__a31o_1
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14127_ clknet_leaf_32_clk _00673_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12388_ _06163_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11339_ sha256cu.m_pad_pars.block_512\[25\]\[2\] _05140_ _05141_ sha256cu.m_pad_pars.block_512\[29\]\[2\]
+ _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__a221o_1
X_14058_ clknet_leaf_39_clk _00604_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13009_ _06494_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__clkbuf_1
X_06880_ sha256cu.msg_scheduler.temp_case _01567_ sha256cu.iter_processing.padding_done
+ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08550_ _03120_ _03122_ _03129_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__a21oi_1
X_07501_ sha256cu.m_out_digest.a_in\[16\] VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__clkbuf_4
X_08481_ sha256cu.m_out_digest.e_in\[22\] _03081_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__xnor2_4
XFILLER_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07432_ _02032_ _02060_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09102_ _02599_ _03587_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__xor2_1
X_07363_ _01994_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__buf_6
XFILLER_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07294_ sha256cu.m_pad_pars.add_out0\[6\] _01937_ sha256cu.m_pad_pars.add_out3\[6\]
+ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__o21a_1
X_09033_ _03520_ _03521_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__and2_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09935_ sha256cu.msg_scheduler.mreg_0\[6\] _04195_ _04199_ _04198_ VGND VGND VPWR
+ VPWR _00466_ sky130_fd_sc_hd__o211a_1
XFILLER_120_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09866_ sha256cu.msg_scheduler.mreg_12\[18\] _04153_ _04156_ _04157_ VGND VGND VPWR
+ VPWR _00433_ sky130_fd_sc_hd__o211a_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08817_ _03313_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ sha256cu.msg_scheduler.mreg_14\[21\] _04106_ VGND VGND VPWR VPWR _04118_
+ sky130_fd_sc_hd__or2_1
XFILLER_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_216 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _03245_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__nand2_1
XANTENNA_205 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08679_ sha256cu.m_out_digest.d_in\[21\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[21\]
+ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__a22o_1
XFILLER_54_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_227 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10710_ sha256cu.msg_scheduler.mreg_10\[19\] _04633_ _04641_ _04636_ VGND VGND VPWR
+ VPWR _00799_ sky130_fd_sc_hd__o211a_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ sha256cu.msg_scheduler.mreg_14\[23\] _05518_ VGND VGND VPWR VPWR _05519_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10641_ sha256cu.msg_scheduler.mreg_9\[21\] _04594_ _04602_ _04597_ VGND VGND VPWR
+ VPWR _00769_ sky130_fd_sc_hd__o211a_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10572_ sha256cu.msg_scheduler.mreg_9\[24\] _04561_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__or2_1
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13360_ _06680_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12311_ _06075_ _06092_ _06113_ _06091_ _06111_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__a221o_1
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13291_ sha256cu.m_pad_pars.block_512\[55\]\[0\] _06644_ VGND VGND VPWR VPWR _06645_
+ sky130_fd_sc_hd__and2_1
X_12242_ _06046_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__nor2_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12173_ _05979_ _05980_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__nand2_1
XFILLER_110_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11124_ sha256cu.m_pad_pars.m_size\[8\] sha256cu.m_pad_pars.block_512\[62\]\[0\]
+ _01919_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__mux2_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11055_ _04755_ _04798_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__and3_1
XFILLER_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10006_ sha256cu.msg_scheduler.mreg_1\[5\] _04234_ _04239_ _04237_ VGND VGND VPWR
+ VPWR _00497_ sky130_fd_sc_hd__o211a_1
XFILLER_103_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14814_ clknet_leaf_117_clk _01328_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11957_ sha256cu.iter_processing.w\[15\] _05666_ _05774_ _05640_ VGND VGND VPWR VPWR
+ _00913_ sky130_fd_sc_hd__o211a_1
X_14745_ clknet_leaf_126_clk _01259_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10908_ _04701_ _04768_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__nor2_2
X_11888_ _05708_ _05706_ _05465_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14676_ clknet_leaf_124_clk _01190_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13627_ clknet_leaf_67_clk _00173_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10839_ sha256cu.msg_scheduler.counter_iteration\[6\] _04185_ _04717_ VGND VGND VPWR
+ VPWR _00852_ sky130_fd_sc_hd__o21a_1
X_13558_ clknet_leaf_65_clk _00104_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_9_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12509_ _06227_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13489_ _06757_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07981_ sha256cu.m_out_digest.g_in\[16\] sha256cu.m_out_digest.f_in\[16\] sha256cu.m_out_digest.e_in\[16\]
+ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__mux2_2
X_09720_ sha256cu.iter_processing.w\[20\] _04067_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__or2_1
X_06932_ _01606_ _01588_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__nand2_1
XFILLER_28_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09651_ sha256cu.m_out_digest.h_in\[15\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[15\]
+ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__o22a_1
X_06863_ _01560_ sha256cu.hashing_done VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__and2b_1
X_09582_ sha256cu.m_out_digest.f_in\[22\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[22\]
+ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__a22o_1
X_08602_ sha256cu.m_out_digest.b_in\[20\] _03179_ _03178_ _02273_ VGND VGND VPWR VPWR
+ _00147_ sky130_fd_sc_hd__a22o_1
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06794_ net213 net216 net215 net218 VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__or4_2
X_08533_ _03114_ _03092_ _03131_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__nand3_1
XFILLER_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08464_ _03064_ _03065_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__nand2_1
X_07415_ sha256cu.m_out_digest.b_in\[1\] sha256cu.m_out_digest.a_in\[1\] sha256cu.m_out_digest.c_in\[1\]
+ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__a21o_1
X_08395_ _02272_ _02997_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07346_ _01986_ _01970_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__nor2_4
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09016_ _03491_ _03492_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__nand2_1
X_07277_ _01927_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09918_ _01567_ sha256cu.iter_processing.padding_done VGND VGND VPWR VPWR _04190_
+ sky130_fd_sc_hd__and2b_1
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09849_ sha256cu.msg_scheduler.mreg_13\[11\] _04147_ VGND VGND VPWR VPWR _04148_
+ sky130_fd_sc_hd__or2_1
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12860_ sha256cu.m_pad_pars.block_512\[29\]\[7\] _05250_ _06351_ VGND VGND VPWR VPWR
+ _06415_ sky130_fd_sc_hd__mux2_1
XFILLER_37_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _05605_ _05610_ _05633_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a21o_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ clknet_leaf_105_clk _01044_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12791_ _06378_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__clkbuf_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ sha256cu.data_in_padd\[6\] _05448_ _05568_ _05463_ VGND VGND VPWR VPWR _05569_
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11673_ _05500_ _05501_ _05433_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__a21oi_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ clknet_leaf_121_clk _00975_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10624_ sha256cu.msg_scheduler.mreg_9\[14\] _04581_ _04592_ _04584_ VGND VGND VPWR
+ VPWR _00762_ sky130_fd_sc_hd__o211a_1
X_14392_ clknet_leaf_47_clk _00906_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[8\]
+ sky130_fd_sc_hd__dfxtp_4
X_13412_ _06707_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13343_ sha256cu.m_pad_pars.block_512\[58\]\[1\] _06671_ VGND VGND VPWR VPWR _06672_
+ sky130_fd_sc_hd__and2_1
XFILLER_10_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10555_ sha256cu.msg_scheduler.mreg_9\[17\] _04548_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__or2_1
X_10486_ _04447_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__buf_2
X_13274_ sha256cu.m_pad_pars.block_512\[54\]\[0\] _06635_ VGND VGND VPWR VPWR _06636_
+ sky130_fd_sc_hd__and2_1
X_12225_ sha256cu.data_in_padd\[26\] _05667_ _06031_ _05445_ VGND VGND VPWR VPWR _06032_
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12156_ _05931_ _05953_ _05955_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11107_ sha256cu.m_pad_pars.add_out2\[4\] sha256cu.m_pad_pars.add_out2\[5\] VGND
+ VGND VPWR VPWR _04966_ sky130_fd_sc_hd__or2b_1
XFILLER_1_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12087_ sha256cu.msg_scheduler.mreg_1\[28\] _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11038_ sha256cu.m_pad_pars.block_512\[31\]\[6\] _04811_ _04828_ sha256cu.m_pad_pars.block_512\[23\]\[6\]
+ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__a22o_1
XFILLER_77_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12989_ sha256cu.m_pad_pars.block_512\[37\]\[3\] _06480_ VGND VGND VPWR VPWR _06484_
+ sky130_fd_sc_hd__and2_1
X_14728_ clknet_leaf_7_clk _01242_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14659_ clknet_leaf_98_clk _01173_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_08180_ _02750_ _02748_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__and2b_1
X_07200_ _01679_ _01860_ _01861_ _01864_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__a31oi_1
XFILLER_146_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07131_ _01593_ _01648_ _01659_ _01804_ _01596_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__a311o_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07062_ _01667_ _01643_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__or2_1
XFILLER_133_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07964_ _02536_ _02534_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__and2b_1
X_07895_ _02482_ _02483_ _02509_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__a21oi_1
X_09703_ sha256cu.msg_scheduler.mreg_14\[12\] _04060_ _04063_ _04064_ VGND VGND VPWR
+ VPWR _00363_ sky130_fd_sc_hd__o211a_1
XFILLER_67_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06915_ _01573_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__buf_4
X_09634_ sha256cu.m_out_digest.h_in\[1\] _04037_ _04036_ sha256cu.m_out_digest.g_in\[1\]
+ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__a22o_1
X_06846_ net248 net251 net250 net253 VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__or4_1
XFILLER_83_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06777_ net201 net234 net223 net256 VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__or4_2
X_09565_ sha256cu.m_out_digest.f_in\[7\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[7\]
+ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__o22a_1
XFILLER_83_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08516_ _02273_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__xnor2_2
X_09496_ _03075_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08447_ _03046_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__xor2_1
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08378_ _02943_ _02959_ _02980_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__or3b_1
XFILLER_149_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07329_ _01564_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__buf_8
X_10340_ sha256cu.msg_scheduler.mreg_5\[20\] _04421_ _04430_ _04424_ VGND VGND VPWR
+ VPWR _00640_ sky130_fd_sc_hd__o211a_1
XFILLER_125_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10271_ sha256cu.msg_scheduler.mreg_4\[23\] _04380_ _04390_ _04383_ VGND VGND VPWR
+ VPWR _00611_ sky130_fd_sc_hd__o211a_1
XFILLER_105_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12010_ sha256cu.msg_scheduler.mreg_1\[25\] _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13961_ clknet_leaf_58_clk _00507_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12912_ sha256cu.m_pad_pars.block_512\[32\]\[7\] _05394_ _06442_ VGND VGND VPWR VPWR
+ _06443_ sky130_fd_sc_hd__mux2_1
XFILLER_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13892_ clknet_leaf_24_clk _00438_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12843_ sha256cu.m_pad_pars.block_512\[28\]\[7\] _05388_ _06351_ VGND VGND VPWR VPWR
+ _06406_ sky130_fd_sc_hd__mux2_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12774_ _06369_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11725_ _05550_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__nand2_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14513_ clknet_leaf_2_clk _01027_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ clknet_leaf_11_clk _00958_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11656_ sha256cu.msg_scheduler.mreg_9\[3\] sha256cu.msg_scheduler.mreg_0\[3\] VGND
+ VGND VPWR VPWR _05486_ sky130_fd_sc_hd__or2_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10607_ sha256cu.msg_scheduler.mreg_10\[7\] _04574_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__or2_1
X_14375_ clknet_leaf_109_clk _00889_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11587_ _04786_ _05275_ sha256cu.m_pad_pars.block_512\[8\]\[7\] VGND VGND VPWR VPWR
+ _05423_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10538_ sha256cu.msg_scheduler.mreg_8\[9\] _04540_ _04542_ _04543_ VGND VGND VPWR
+ VPWR _00725_ sky130_fd_sc_hd__o211a_1
XFILLER_6_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13326_ sha256cu.m_pad_pars.block_512\[57\]\[1\] _06660_ VGND VGND VPWR VPWR _06663_
+ sky130_fd_sc_hd__and2_1
XFILLER_115_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13257_ sha256cu.m_pad_pars.block_512\[53\]\[0\] _06626_ VGND VGND VPWR VPWR _06627_
+ sky130_fd_sc_hd__and2_1
X_10469_ sha256cu.msg_scheduler.mreg_8\[12\] _04494_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__or2_1
X_12208_ _06012_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__xor2_1
XFILLER_142_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13188_ _05269_ _06589_ _01972_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__o21ai_4
X_12139_ _05946_ _05947_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__and2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07680_ sha256cu.m_out_digest.e_in\[19\] _02301_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__xnor2_4
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09350_ _03826_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__and2_1
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09281_ _02777_ _03729_ _03730_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__a21boi_1
X_08301_ _02889_ _02890_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__a21oi_1
X_08232_ _02761_ _02801_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__or2_1
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08163_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__inv_2
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08094_ sha256cu.iter_processing.w\[18\] _02672_ _02704_ VGND VGND VPWR VPWR _02705_
+ sky130_fd_sc_hd__a21o_1
X_07114_ _01620_ _01780_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__or2_1
X_07045_ _00454_ _01727_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__nor2_1
XFILLER_142_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08996_ _03481_ _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__nor2_1
XFILLER_114_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07947_ _02560_ _02561_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__xnor2_2
XFILLER_88_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07878_ _02161_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__xnor2_2
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06829_ _01523_ _01524_ _01525_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__or4_1
X_09617_ sha256cu.m_out_digest.g_in\[19\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[19\]
+ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__a22o_1
XFILLER_44_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09548_ _03992_ _03996_ _03990_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__o21a_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09479_ _03951_ _03952_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__nand2_1
X_11510_ sha256cu.m_pad_pars.block_512\[20\]\[3\] _05294_ _05285_ sha256cu.m_pad_pars.block_512\[16\]\[3\]
+ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__a22o_1
XFILLER_12_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12490_ _06217_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11441_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__inv_1
X_14160_ clknet_leaf_31_clk _00706_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11372_ sha256cu.m_pad_pars.block_512\[49\]\[5\] _05151_ _05158_ sha256cu.m_pad_pars.block_512\[21\]\[5\]
+ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__a221o_1
X_10323_ sha256cu.msg_scheduler.mreg_5\[13\] _04407_ _04420_ _04410_ VGND VGND VPWR
+ VPWR _00633_ sky130_fd_sc_hd__o211a_1
X_13111_ sha256cu.m_pad_pars.block_512\[44\]\[4\] _06544_ VGND VGND VPWR VPWR _06549_
+ sky130_fd_sc_hd__and2_1
X_14091_ clknet_leaf_37_clk _00637_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10254_ sha256cu.msg_scheduler.mreg_5\[16\] _04374_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__or2_1
XFILLER_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13042_ sha256cu.m_pad_pars.block_512\[40\]\[4\] _06507_ VGND VGND VPWR VPWR _06512_
+ sky130_fd_sc_hd__and2_1
X_10185_ sha256cu.msg_scheduler.mreg_4\[18\] _04335_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__or2_1
XFILLER_132_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13944_ clknet_leaf_43_clk _00490_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13875_ clknet_leaf_20_clk _00421_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12826_ sha256cu.m_pad_pars.block_512\[27\]\[7\] _04945_ _06351_ VGND VGND VPWR VPWR
+ _06397_ sky130_fd_sc_hd__mux2_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12757_ _06360_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__clkbuf_1
X_11708_ _05508_ _05512_ _05509_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__a21boi_1
X_12688_ _06323_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_1
X_11639_ _05468_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__nand2_1
X_14427_ clknet_leaf_100_clk _00941_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14358_ clknet_leaf_110_clk _00872_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13309_ sha256cu.m_pad_pars.block_512\[56\]\[1\] _01924_ VGND VGND VPWR VPWR _06654_
+ sky130_fd_sc_hd__and2_1
XFILLER_131_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14289_ clknet_leaf_25_clk _00835_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08850_ sha256cu.iter_processing.w\[7\] _02264_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__nand2_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07801_ _02083_ _02419_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__xnor2_2
XFILLER_97_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08781_ _03276_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__xnor2_1
X_07732_ _02342_ _02352_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__xor2_1
XFILLER_37_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07663_ _02243_ _02241_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__and2b_1
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09402_ sha256cu.iter_processing.w\[26\] _02971_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__nor2_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07594_ _01913_ _02218_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__or2_1
XFILLER_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09333_ sha256cu.m_out_digest.e_in\[23\] _02439_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__or2_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_126_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_34_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09264_ _03701_ _03708_ _03743_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__or3_1
XFILLER_21_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09195_ sha256cu.iter_processing.w\[19\] _02708_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__nand2_1
X_08215_ _02821_ _02822_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__nor2_1
X_08146_ _02737_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__xnor2_2
X_08077_ _02668_ _02687_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__nor2_1
XFILLER_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07028_ _01655_ _01689_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__nor2_1
XFILLER_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08979_ _03450_ _03451_ _03468_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11990_ _05803_ _05804_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__and2_1
XFILLER_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10941_ _04748_ _04776_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__or2_2
X_13660_ clknet_leaf_68_clk _00206_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12611_ sha256cu.m_pad_pars.block_512\[15\]\[2\] _06280_ VGND VGND VPWR VPWR _06283_
+ sky130_fd_sc_hd__and2_1
X_10872_ _02002_ _01960_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__nor2_1
X_13591_ clknet_leaf_63_clk _00137_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_117_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12542_ sha256cu.m_pad_pars.block_512\[11\]\[3\] _06241_ VGND VGND VPWR VPWR _06245_
+ sky130_fd_sc_hd__and2_1
X_12473_ _06208_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14212_ clknet_leaf_28_clk _00758_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11424_ sha256cu.m_pad_pars.block_512\[61\]\[7\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[7\]
+ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__a22o_1
XFILLER_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_35_clk _00689_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11355_ sha256cu.m_pad_pars.block_512\[13\]\[4\] _05128_ _05147_ sha256cu.m_pad_pars.block_512\[33\]\[4\]
+ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a221o_1
XFILLER_153_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10306_ sha256cu.msg_scheduler.mreg_6\[6\] _04401_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__or2_1
X_14074_ clknet_leaf_44_clk _00620_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11286_ _04807_ _05004_ _05136_ _04805_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__o22a_1
XFILLER_152_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10237_ sha256cu.msg_scheduler.mreg_4\[8\] _04367_ _04371_ _04370_ VGND VGND VPWR
+ VPWR _00596_ sky130_fd_sc_hd__o211a_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13025_ sha256cu.m_pad_pars.block_512\[39\]\[4\] _06498_ VGND VGND VPWR VPWR _06503_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10168_ sha256cu.msg_scheduler.mreg_3\[10\] _04328_ _04332_ _04331_ VGND VGND VPWR
+ VPWR _00566_ sky130_fd_sc_hd__o211a_1
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10099_ sha256cu.msg_scheduler.mreg_3\[13\] _04282_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__or2_1
XFILLER_82_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13927_ clknet_leaf_43_clk _00473_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13858_ clknet_leaf_23_clk _00404_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13789_ clknet_leaf_68_clk _00335_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12809_ sha256cu.m_pad_pars.block_512\[26\]\[7\] _05083_ _06351_ VGND VGND VPWR VPWR
+ _06388_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_16_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08000_ _02558_ _02577_ _02613_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__a21o_1
XFILLER_144_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09951_ _04166_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08902_ _03368_ _03385_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__nand2_1
XFILLER_131_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09882_ _04043_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _03316_ _03317_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__o21ai_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _03255_ _03257_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__nor2_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ sha256cu.m_out_digest.b_in\[9\] sha256cu.m_out_digest.a_in\[9\] VGND VGND
+ VPWR VPWR _02336_ sky130_fd_sc_hd__or2_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08695_ _03195_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nand2_1
XANTENNA_409 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07646_ sha256cu.m_out_digest.e_in\[13\] sha256cu.m_out_digest.e_in\[0\] VGND VGND
+ VPWR VPWR _02269_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07577_ _02197_ _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09316_ sha256cu.iter_processing.w\[23\] _02859_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__or2_1
XFILLER_139_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09247_ _03713_ _03714_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__nand2_1
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09178_ _03630_ _03642_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__a21oi_1
X_08129_ sha256cu.m_out_digest.b_in\[20\] _02273_ _02738_ VGND VGND VPWR VPWR _02739_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11140_ _04997_ _04998_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__nor2_2
XFILLER_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 hash[190] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
X_11071_ sha256cu.m_pad_pars.block_512\[59\]\[7\] _04829_ _04906_ _04916_ _04930_
+ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__a2111o_1
Xinput123 hash[20] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput145 hash[22] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlymetal6s2s_1
X_10022_ sha256cu.msg_scheduler.mreg_1\[12\] _04247_ _04248_ _04237_ VGND VGND VPWR
+ VPWR _00504_ sky130_fd_sc_hd__o211a_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput134 hash[21] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xinput112 hash[1] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 hash[24] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
Xinput156 hash[23] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
X_14830_ clknet_leaf_113_clk _01344_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput178 hash[29] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput189 hash[39] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_2
XFILLER_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11973_ _05788_ _05789_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__nand2_1
X_14761_ clknet_leaf_16_clk _01275_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13712_ clknet_leaf_66_clk _00258_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10924_ _04743_ sha256cu.m_pad_pars.add_512_block\[4\] VGND VGND VPWR VPWR _04791_
+ sky130_fd_sc_hd__or2_4
X_14692_ clknet_leaf_103_clk _01206_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13643_ clknet_leaf_74_clk _00189_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10855_ sha256cu.m_pad_pars.add_out3\[2\] _01963_ _01966_ VGND VGND VPWR VPWR _04729_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_32_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13574_ clknet_leaf_85_clk _00120_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[25\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_13_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10786_ sha256cu.msg_scheduler.mreg_12\[21\] _04679_ VGND VGND VPWR VPWR _04684_
+ sky130_fd_sc_hd__or2_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ sha256cu.m_pad_pars.block_512\[10\]\[3\] _06232_ VGND VGND VPWR VPWR _06236_
+ sky130_fd_sc_hd__and2_1
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12456_ _06199_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12387_ sha256cu.m_pad_pars.block_512\[2\]\[2\] _06160_ VGND VGND VPWR VPWR _06163_
+ sky130_fd_sc_hd__and2_1
X_11407_ _01977_ _01985_ _05250_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__and3_1
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14126_ clknet_leaf_32_clk _00672_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11338_ sha256cu.m_pad_pars.block_512\[5\]\[2\] _05160_ _05161_ sha256cu.m_pad_pars.block_512\[53\]\[2\]
+ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a221o_1
XFILLER_140_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14057_ clknet_leaf_40_clk _00603_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11269_ _04917_ _04993_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__o21ai_1
X_13008_ sha256cu.m_pad_pars.block_512\[38\]\[4\] _06489_ VGND VGND VPWR VPWR _06494_
+ sky130_fd_sc_hd__and2_1
XFILLER_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07500_ _02126_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__inv_2
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14959_ clknet_leaf_95_clk _01473_ VGND VGND VPWR VPWR sha256cu.temp_case sky130_fd_sc_hd__dfxtp_1
X_08480_ sha256cu.m_out_digest.e_in\[8\] sha256cu.m_out_digest.e_in\[3\] VGND VGND
+ VPWR VPWR _03081_ sky130_fd_sc_hd__xnor2_4
XFILLER_35_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07431_ _02049_ _02059_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__xor2_1
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07362_ _01976_ _01998_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__nand2_1
X_09101_ _03585_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nand2_1
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07293_ _01935_ _01936_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__nand2_2
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09032_ _03506_ _03486_ _03519_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__or3_1
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09934_ sha256cu.msg_scheduler.mreg_1\[6\] _04174_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__or2_1
X_09865_ _04116_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__buf_2
XFILLER_86_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _02002_ _03312_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__or2_1
XFILLER_100_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09796_ sha256cu.msg_scheduler.mreg_13\[20\] _04112_ _04115_ _04117_ VGND VGND VPWR
+ VPWR _00403_ sky130_fd_sc_hd__o211a_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ sha256cu.m_out_digest.h_in\[3\] sha256cu.m_out_digest.d_in\[3\] VGND VGND
+ VPWR VPWR _03246_ sky130_fd_sc_hd__nand2_1
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_206 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_217 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_239 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ sha256cu.m_out_digest.d_in\[20\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[20\]
+ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__a22o_1
XANTENNA_228 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07629_ _02178_ _02180_ _02186_ _02214_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__o22a_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10640_ sha256cu.msg_scheduler.mreg_10\[21\] _04601_ VGND VGND VPWR VPWR _04602_
+ sky130_fd_sc_hd__or2_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10571_ sha256cu.msg_scheduler.mreg_8\[23\] _04554_ _04562_ _04557_ VGND VGND VPWR
+ VPWR _00739_ sky130_fd_sc_hd__o211a_1
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12310_ _06072_ _06090_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__or2_1
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13290_ _01986_ _04832_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__or2_2
X_12241_ _06017_ _06021_ _06044_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12172_ _05979_ _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__or2_1
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11123_ _04725_ sha256cu.m_pad_pars.add_out2\[4\] _04958_ VGND VGND VPWR VPWR _04982_
+ sky130_fd_sc_hd__and3_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11054_ _04753_ _04913_ _04802_ sha256cu.m_pad_pars.block_512\[43\]\[7\] VGND VGND
+ VPWR VPWR _04914_ sky130_fd_sc_hd__o22a_1
X_10005_ sha256cu.msg_scheduler.mreg_2\[5\] _04228_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__or2_1
XFILLER_92_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14813_ clknet_leaf_119_clk _01327_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11956_ sha256cu.data_in_padd\[15\] _05667_ _05773_ _05445_ VGND VGND VPWR VPWR _05774_
+ sky130_fd_sc_hd__a211o_1
X_14744_ clknet_leaf_120_clk _01258_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10907_ _04766_ _04767_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__and3_2
XFILLER_32_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11887_ _05658_ _05662_ _05682_ _05681_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__a31o_1
X_14675_ clknet_leaf_1_clk _01189_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13626_ clknet_leaf_67_clk _00172_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10838_ sha256cu.msg_scheduler.counter_iteration\[6\] _04185_ _04177_ VGND VGND VPWR
+ VPWR _04717_ sky130_fd_sc_hd__a21oi_1
XFILLER_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13557_ clknet_leaf_61_clk _00103_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[8\]
+ sky130_fd_sc_hd__dfxtp_4
X_10769_ _01994_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__buf_2
XFILLER_146_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12508_ sha256cu.m_pad_pars.block_512\[9\]\[3\] _06223_ VGND VGND VPWR VPWR _06227_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13488_ _06730_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__and2_1
X_12439_ _06190_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ clknet_leaf_36_clk _00655_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07980_ sha256cu.m_out_digest.b_in\[16\] _02128_ _02593_ VGND VGND VPWR VPWR _02594_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_86_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06931_ _00454_ _01608_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__nor2_2
X_09650_ sha256cu.m_out_digest.h_in\[14\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[14\]
+ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__o22a_1
XFILLER_95_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08601_ _02923_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__buf_6
X_06862_ _01503_ _01517_ _01538_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__nor4_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06793_ _01487_ _01488_ _01489_ _01490_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__or4_2
X_09581_ sha256cu.m_out_digest.f_in\[21\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[21\]
+ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__a22o_1
X_08532_ _03114_ _03092_ _03131_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__a21o_1
X_08463_ _03038_ _03039_ _03063_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__or3b_1
X_07414_ sha256cu.m_out_digest.b_in\[1\] sha256cu.m_out_digest.a_in\[1\] VGND VGND
+ VPWR VPWR _02043_ sky130_fd_sc_hd__or2_1
XFILLER_51_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08394_ _02162_ sha256cu.m_out_digest.a_in\[8\] VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07345_ _01911_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__buf_4
XFILLER_148_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
X_07276_ sha256cu.m_pad_pars.block_512\[63\]\[2\] _01924_ VGND VGND VPWR VPWR _01927_
+ sky130_fd_sc_hd__and2_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09015_ sha256cu.m_out_digest.e_in\[12\] _02732_ _03503_ _03504_ _02258_ VGND VGND
+ VPWR VPWR _00235_ sky130_fd_sc_hd__a221o_1
XFILLER_152_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09917_ sha256cu.msg_scheduler.counter_iteration\[6\] _01574_ _04189_ _04171_ VGND
+ VGND VPWR VPWR _00458_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_97_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
X_09848_ _04133_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__clkbuf_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09779_ sha256cu.msg_scheduler.mreg_13\[13\] _04099_ _04107_ _04103_ VGND VGND VPWR
+ VPWR _00396_ sky130_fd_sc_hd__o211a_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _05605_ _05610_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__nand3_1
XFILLER_74_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12790_ sha256cu.m_pad_pars.block_512\[25\]\[6\] _06371_ VGND VGND VPWR VPWR _06378_
+ sky130_fd_sc_hd__and2_1
XFILLER_27_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _05465_ _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__nor2_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _05500_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__or2_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14460_ clknet_leaf_126_clk _00974_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10623_ sha256cu.msg_scheduler.mreg_10\[14\] _04588_ VGND VGND VPWR VPWR _04592_
+ sky130_fd_sc_hd__or2_1
X_14391_ clknet_leaf_15_clk _00905_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[7\]
+ sky130_fd_sc_hd__dfxtp_4
X_13411_ sha256cu.m_pad_pars.block_512\[62\]\[2\] _01928_ VGND VGND VPWR VPWR _06707_
+ sky130_fd_sc_hd__and2_1
XFILLER_128_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10554_ sha256cu.msg_scheduler.mreg_8\[16\] _04540_ _04552_ _04543_ VGND VGND VPWR
+ VPWR _00732_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_21_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13342_ _01923_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10485_ sha256cu.msg_scheduler.mreg_7\[19\] _04500_ _04512_ _04503_ VGND VGND VPWR
+ VPWR _00703_ sky130_fd_sc_hd__o211a_1
XFILLER_136_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13273_ _04979_ _04980_ _01912_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__a21o_2
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12224_ _06026_ _06029_ _06030_ _05465_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__a211oi_1
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12155_ _05933_ _05936_ _05956_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__or3b_1
XFILLER_45_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11106_ sha256cu.m_pad_pars.block_512\[10\]\[0\] _04963_ _04964_ sha256cu.m_pad_pars.block_512\[26\]\[0\]
+ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__a22o_1
X_12086_ sha256cu.msg_scheduler.mreg_1\[24\] sha256cu.msg_scheduler.mreg_1\[7\] VGND
+ VGND VPWR VPWR _05898_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_88_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_65_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11037_ sha256cu.m_pad_pars.block_512\[27\]\[6\] _04757_ _04804_ sha256cu.m_pad_pars.block_512\[43\]\[6\]
+ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__a22o_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12988_ _06483_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__clkbuf_1
X_11939_ _05755_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__nand2_1
X_14727_ clknet_leaf_12_clk _01241_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14658_ clknet_leaf_96_clk _01172_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13609_ clknet_leaf_78_clk _00155_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
X_14589_ clknet_leaf_117_clk _01103_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_07130_ _01632_ _01659_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__nor2_1
XFILLER_9_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07061_ _00455_ _01670_ _01675_ _00456_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__a211o_1
XFILLER_99_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07963_ _02558_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__xnor2_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
X_07894_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__inv_2
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09702_ _01973_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__buf_2
X_06914_ _01577_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__nand2_4
XFILLER_28_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09633_ sha256cu.m_out_digest.h_in\[0\] _04035_ _04038_ sha256cu.m_out_digest.g_in\[0\]
+ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__o22a_1
X_06845_ _01539_ _01540_ _01541_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__or4_1
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09564_ _02515_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__buf_4
XFILLER_56_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08515_ sha256cu.m_out_digest.a_in\[11\] sha256cu.m_out_digest.a_in\[0\] VGND VGND
+ VPWR VPWR _03115_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06776_ _01474_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__clkbuf_1
X_09495_ _03966_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__nand2_1
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08446_ sha256cu.m_out_digest.h_in\[27\] _02998_ _03047_ VGND VGND VPWR VPWR _03048_
+ sky130_fd_sc_hd__a21bo_1
X_08377_ _02943_ _02959_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__o21ba_1
XFILLER_11_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07328_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__buf_4
XFILLER_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07259_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__buf_6
X_10270_ sha256cu.msg_scheduler.mreg_5\[23\] _04387_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__or2_1
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13960_ clknet_leaf_59_clk _00506_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12911_ _01964_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__buf_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13891_ clknet_leaf_24_clk _00437_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12842_ _06405_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__clkbuf_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ sha256cu.m_pad_pars.block_512\[24\]\[6\] _06362_ VGND VGND VPWR VPWR _06369_
+ sky130_fd_sc_hd__and2_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11724_ sha256cu.msg_scheduler.mreg_9\[6\] sha256cu.msg_scheduler.mreg_0\[6\] VGND
+ VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nand2_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ clknet_leaf_2_clk _01026_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11655_ sha256cu.msg_scheduler.mreg_9\[3\] sha256cu.msg_scheduler.mreg_0\[3\] VGND
+ VGND VPWR VPWR _05485_ sky130_fd_sc_hd__nand2_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14443_ clknet_leaf_9_clk _00957_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10606_ sha256cu.msg_scheduler.mreg_9\[6\] _04581_ _04582_ _04570_ VGND VGND VPWR
+ VPWR _00754_ sky130_fd_sc_hd__o211a_1
X_14374_ clknet_leaf_110_clk _00888_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11586_ _01920_ _05419_ _05421_ _05287_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__a22o_1
X_10537_ _04529_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__buf_2
XFILLER_6_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13325_ _06662_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_1
X_10468_ sha256cu.msg_scheduler.mreg_7\[11\] _04500_ _04502_ _04503_ VGND VGND VPWR
+ VPWR _00695_ sky130_fd_sc_hd__o211a_1
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13256_ _02111_ _01950_ _04705_ _05159_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__or4_4
X_12207_ sha256cu.msg_scheduler.mreg_1\[29\] _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10399_ sha256cu.msg_scheduler.mreg_6\[13\] _04461_ _04463_ _04464_ VGND VGND VPWR
+ VPWR _00665_ sky130_fd_sc_hd__o211a_1
XFILLER_124_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13187_ _01952_ _05136_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__nor2_1
X_12138_ _05946_ _05947_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__nor2_1
XFILLER_96_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12069_ _05854_ _05856_ _05852_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_77_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09280_ _02811_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__xor2_1
X_08300_ _02900_ _02905_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__xnor2_1
X_08231_ _02837_ _02838_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__or2_1
XFILLER_21_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08162_ sha256cu.iter_processing.w\[20\] _02741_ _02770_ VGND VGND VPWR VPWR _02771_
+ sky130_fd_sc_hd__a21o_1
XFILLER_109_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08093_ _02670_ _02671_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__and2b_1
X_07113_ _01701_ _01704_ _01705_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__a21o_1
X_07044_ _01580_ _01590_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__nand2_1
XFILLER_115_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08995_ sha256cu.K\[12\] _03484_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07946_ sha256cu.m_out_digest.g_in\[15\] sha256cu.m_out_digest.f_in\[15\] sha256cu.m_out_digest.e_in\[15\]
+ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__mux2_2
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07877_ _02084_ sha256cu.m_out_digest.a_in\[3\] VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06828_ net72 net75 net74 net77 VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__or4_2
X_09616_ sha256cu.m_out_digest.g_in\[18\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[18\]
+ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__a22o_1
X_09547_ _04000_ _04001_ _03998_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09478_ _03948_ _03950_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__or2_1
XFILLER_24_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08429_ _02069_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11440_ _01944_ _04699_ _04777_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__a31o_1
XFILLER_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11371_ sha256cu.m_pad_pars.block_512\[5\]\[5\] _05160_ _05161_ sha256cu.m_pad_pars.block_512\[53\]\[5\]
+ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__a221o_1
X_14090_ clknet_leaf_33_clk _00636_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10322_ sha256cu.msg_scheduler.mreg_6\[13\] _04415_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__or2_1
XFILLER_3_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13110_ _06548_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_1
X_13041_ _06511_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__clkbuf_1
X_10253_ _04314_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__buf_2
XFILLER_79_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10184_ _04314_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__buf_2
XFILLER_79_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13943_ clknet_leaf_46_clk _00489_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_13874_ clknet_leaf_18_clk _00420_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12825_ _06396_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__clkbuf_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ sha256cu.m_pad_pars.block_512\[23\]\[6\] _06353_ VGND VGND VPWR VPWR _06360_
+ sky130_fd_sc_hd__and2_1
X_11707_ _05532_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__xor2_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ sha256cu.m_pad_pars.block_512\[19\]\[6\] _06316_ VGND VGND VPWR VPWR _06323_
+ sky130_fd_sc_hd__and2_1
X_11638_ sha256cu.msg_scheduler.mreg_9\[2\] sha256cu.msg_scheduler.mreg_0\[2\] VGND
+ VGND VPWR VPWR _05469_ sky130_fd_sc_hd__or2_1
X_14426_ clknet_leaf_118_clk _00940_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14357_ clknet_leaf_110_clk _00871_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13308_ _06653_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
X_11569_ _04908_ _04924_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14288_ clknet_leaf_25_clk _00834_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13239_ _06270_ _05308_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__nand2_2
X_08780_ _03244_ _03250_ _03277_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__o21a_1
X_07800_ _02027_ sha256cu.m_out_digest.a_in\[1\] VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__xnor2_1
X_07731_ _02349_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07662_ _02261_ _02284_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__xnor2_2
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07593_ sha256cu.m_out_digest.a_in\[5\] _02037_ _02017_ _02217_ VGND VGND VPWR VPWR
+ _02218_ sky130_fd_sc_hd__a22o_1
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09401_ _03875_ _03876_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__nand2_1
XFILLER_111_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09332_ _03777_ _03784_ _03809_ _02629_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__a31o_1
XFILLER_52_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09263_ _03701_ _03708_ _03743_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09194_ sha256cu.iter_processing.w\[19\] _02708_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__or2_1
X_08214_ sha256cu.iter_processing.w\[22\] _02820_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__and2_1
XFILLER_21_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08145_ _02752_ _02754_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__xnor2_2
XFILLER_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08076_ _02668_ _02687_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__and2_1
XFILLER_1_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07027_ _01710_ _01687_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__nor2_1
XFILLER_130_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08978_ _03450_ _03451_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__and3_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07929_ _02542_ _02544_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__xor2_2
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10940_ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__clkbuf_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12610_ _06282_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__clkbuf_1
X_10871_ sha256cu.m_pad_pars.add_out3\[6\] _04739_ _04740_ VGND VGND VPWR VPWR _00861_
+ sky130_fd_sc_hd__o21ba_1
X_13590_ clknet_leaf_63_clk _00136_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12541_ _06244_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12472_ sha256cu.m_pad_pars.block_512\[7\]\[2\] _06205_ VGND VGND VPWR VPWR _06208_
+ sky130_fd_sc_hd__and2_1
XFILLER_12_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14211_ clknet_leaf_28_clk _00757_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11423_ _05264_ _04913_ _05145_ sha256cu.m_pad_pars.block_512\[33\]\[7\] VGND VGND
+ VPWR VPWR _05267_ sky130_fd_sc_hd__o22a_1
XFILLER_138_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14142_ clknet_leaf_36_clk _00688_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11354_ sha256cu.m_pad_pars.block_512\[45\]\[4\] _05126_ VGND VGND VPWR VPWR _05201_
+ sky130_fd_sc_hd__and2_1
XFILLER_4_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10305_ sha256cu.msg_scheduler.mreg_5\[5\] _04407_ _04409_ _04410_ VGND VGND VPWR
+ VPWR _00625_ sky130_fd_sc_hd__o211a_1
X_14073_ clknet_leaf_44_clk _00619_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11285_ _01942_ _04699_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__nand2_4
X_10236_ sha256cu.msg_scheduler.mreg_5\[8\] _04361_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__or2_1
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13024_ _06502_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10167_ sha256cu.msg_scheduler.mreg_4\[10\] _04322_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__or2_1
XFILLER_121_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10098_ sha256cu.msg_scheduler.mreg_2\[12\] _04288_ _04292_ _04291_ VGND VGND VPWR
+ VPWR _00536_ sky130_fd_sc_hd__o211a_1
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13926_ clknet_leaf_44_clk _00472_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13857_ clknet_leaf_23_clk _00403_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13788_ clknet_leaf_68_clk _00334_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_12808_ _06387_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__clkbuf_1
X_12739_ _06350_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__clkbuf_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14409_ clknet_leaf_77_clk _00923_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[25\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_129_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09950_ sha256cu.msg_scheduler.mreg_0\[13\] _04195_ _04207_ _04198_ VGND VGND VPWR
+ VPWR _00473_ sky130_fd_sc_hd__o211a_1
X_08901_ _03384_ _03382_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__or2b_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09881_ sha256cu.msg_scheduler.mreg_12\[25\] _04153_ _04165_ _04157_ VGND VGND VPWR
+ VPWR _00440_ sky130_fd_sc_hd__o211a_1
XFILLER_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _03321_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__xor2_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ sha256cu.m_out_digest.e_in\[4\] VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__inv_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07714_ sha256cu.iter_processing.w\[8\] _02298_ _02297_ VGND VGND VPWR VPWR _02335_
+ sky130_fd_sc_hd__a21o_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08694_ sha256cu.K\[0\] _03193_ _03194_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__nand3_1
XFILLER_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07645_ sha256cu.iter_processing.w\[7\] _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__xnor2_2
X_07576_ sha256cu.m_out_digest.h_in\[5\] _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09315_ sha256cu.K\[23\] VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__inv_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09246_ _02040_ _03726_ _03727_ _03366_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__o211a_1
XFILLER_21_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09177_ _03659_ _03660_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08128_ sha256cu.m_out_digest.b_in\[20\] _02273_ sha256cu.m_out_digest.c_in\[20\]
+ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__a21o_1
X_08059_ sha256cu.m_out_digest.g_in\[18\] sha256cu.m_out_digest.f_in\[18\] sha256cu.m_out_digest.e_in\[18\]
+ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_150_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11070_ _04821_ _04919_ _04921_ _04929_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__a211o_1
Xinput102 hash[191] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10021_ sha256cu.msg_scheduler.mreg_2\[12\] _04241_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__or2_1
XFILLER_88_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput113 hash[200] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_4
Xinput135 hash[220] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xinput124 hash[210] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_2
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput146 hash[230] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput168 hash[250] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_2
Xinput157 hash[240] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14760_ clknet_leaf_12_clk _01274_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput179 hash[2] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13711_ clknet_leaf_73_clk _00257_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11972_ _05785_ _05787_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__or2_1
XFILLER_71_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10923_ _04784_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__nor2_4
X_14691_ clknet_leaf_103_clk _01205_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13642_ clknet_leaf_82_clk _00188_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10854_ sha256cu.m_pad_pars.add_out3\[2\] _01961_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__and2_1
XFILLER_44_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ clknet_leaf_86_clk _00119_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10785_ sha256cu.msg_scheduler.mreg_11\[20\] _04672_ _04683_ _04675_ VGND VGND VPWR
+ VPWR _00832_ sky130_fd_sc_hd__o211a_1
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _06235_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12455_ sha256cu.m_pad_pars.block_512\[6\]\[2\] _06196_ VGND VGND VPWR VPWR _06199_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12386_ _06162_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__clkbuf_1
X_11406_ _04699_ _04925_ _04973_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__a31o_1
X_14125_ clknet_leaf_32_clk _00671_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11337_ sha256cu.m_pad_pars.block_512\[37\]\[2\] _05165_ _05185_ _05024_ VGND VGND
+ VPWR VPWR _05186_ sky130_fd_sc_hd__a22o_1
XFILLER_113_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14056_ clknet_leaf_40_clk _00602_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11268_ _04801_ _05117_ sha256cu.m_pad_pars.block_512\[34\]\[7\] VGND VGND VPWR VPWR
+ _05120_ sky130_fd_sc_hd__a21o_1
X_10219_ _04281_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__clkbuf_2
X_13007_ _06493_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__clkbuf_1
X_11199_ sha256cu.m_pad_pars.block_512\[42\]\[4\] _05001_ _04989_ sha256cu.m_pad_pars.block_512\[14\]\[4\]
+ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__a22o_1
XFILLER_82_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14958_ clknet_leaf_90_clk _01472_ VGND VGND VPWR VPWR sha256cu.K\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_35_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14889_ clknet_leaf_10_clk _01403_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13909_ clknet_leaf_96_clk _00455_ VGND VGND VPWR VPWR sha256cu.counter_iteration\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_07430_ _02056_ _02058_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07361_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__clkbuf_4
X_09100_ sha256cu.m_out_digest.h_in\[16\] sha256cu.m_out_digest.d_in\[16\] VGND VGND
+ VPWR VPWR _03586_ sky130_fd_sc_hd__nand2_1
XFILLER_148_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09031_ _03506_ _03486_ _03519_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__o21ai_1
X_07292_ sha256cu.m_pad_pars.add_out0\[5\] sha256cu.m_pad_pars.add_out0\[4\] VGND
+ VGND VPWR VPWR _01936_ sky130_fd_sc_hd__nor2_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09933_ sha256cu.msg_scheduler.mreg_0\[5\] _04195_ _04197_ _04198_ VGND VGND VPWR
+ VPWR _00465_ sky130_fd_sc_hd__o211a_1
XFILLER_98_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09864_ sha256cu.msg_scheduler.mreg_13\[18\] _04147_ VGND VGND VPWR VPWR _04156_
+ sky130_fd_sc_hd__or2_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08815_ sha256cu.m_out_digest.e_in\[5\] _02037_ _02017_ _03311_ VGND VGND VPWR VPWR
+ _03312_ sky130_fd_sc_hd__a22o_1
XFILLER_112_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__buf_2
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ sha256cu.m_out_digest.h_in\[3\] sha256cu.m_out_digest.d_in\[3\] VGND VGND
+ VPWR VPWR _03245_ sky130_fd_sc_hd__or2_1
XFILLER_54_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_207 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_218 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ sha256cu.m_out_digest.d_in\[19\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[19\]
+ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__o22a_1
XANTENNA_229 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07628_ _02249_ _02251_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__xnor2_2
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07559_ sha256cu.m_out_digest.a_in\[4\] _02070_ _02183_ _02184_ VGND VGND VPWR VPWR
+ _00099_ sky130_fd_sc_hd__a22o_1
X_10570_ sha256cu.msg_scheduler.mreg_9\[23\] _04561_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__or2_1
X_09229_ _03695_ _03681_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__o21ai_1
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12240_ _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__inv_2
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12171_ _05950_ _05951_ _05948_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11122_ _04978_ _04979_ _04980_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__and3_2
XFILLER_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11053_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__buf_4
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10004_ sha256cu.msg_scheduler.mreg_1\[4\] _04234_ _04238_ _04237_ VGND VGND VPWR
+ VPWR _00496_ sky130_fd_sc_hd__o211a_1
XFILLER_67_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14812_ clknet_leaf_117_clk _01326_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11955_ _05771_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__nor2_1
X_14743_ clknet_leaf_120_clk _01257_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14674_ clknet_leaf_1_clk _01188_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10906_ _04702_ _04769_ _04770_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__o31a_1
X_13625_ clknet_leaf_64_clk _00171_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11886_ _05658_ _05662_ _05682_ _05706_ _05681_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__a311o_2
XFILLER_9_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10837_ _04176_ _04715_ _04716_ sha256cu.iter_processing.padding_done _01984_ VGND
+ VGND VPWR VPWR _00851_ sky130_fd_sc_hd__o221ai_1
X_13556_ clknet_leaf_59_clk _00102_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[7\]
+ sky130_fd_sc_hd__dfxtp_4
X_10768_ sha256cu.msg_scheduler.mreg_12\[13\] _04666_ VGND VGND VPWR VPWR _04674_
+ sky130_fd_sc_hd__or2_1
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12507_ _06226_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
X_13487_ sha256cu.K\[21\] _06713_ _06718_ _00049_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__a22o_1
X_10699_ sha256cu.msg_scheduler.mreg_11\[15\] _04627_ VGND VGND VPWR VPWR _04635_
+ sky130_fd_sc_hd__or2_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12438_ sha256cu.m_pad_pars.block_512\[5\]\[2\] _06187_ VGND VGND VPWR VPWR _06190_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12369_ sha256cu.m_pad_pars.block_512\[1\]\[1\] _06152_ VGND VGND VPWR VPWR _06154_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14108_ clknet_leaf_36_clk _00654_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14039_ clknet_leaf_41_clk _00585_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06930_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06861_ _01543_ _01548_ _01553_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__or4_1
X_08600_ sha256cu.m_out_digest.b_in\[19\] _03031_ _03178_ _02233_ VGND VGND VPWR VPWR
+ _00146_ sky130_fd_sc_hd__a22o_1
XFILLER_67_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06792_ net186 net189 net188 net192 VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__or4_2
XFILLER_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09580_ sha256cu.m_out_digest.f_in\[20\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[20\]
+ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__a22o_1
XFILLER_67_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08531_ _03129_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__or2_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08462_ _03038_ _03039_ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__o21bai_1
X_07413_ sha256cu.iter_processing.w\[0\] _02021_ _02041_ VGND VGND VPWR VPWR _02042_
+ sky130_fd_sc_hd__a21o_1
XFILLER_90_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08393_ sha256cu.K\[27\] VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__inv_2
XFILLER_148_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07344_ sha256cu.m_pad_pars.add_out1\[5\] sha256cu.m_pad_pars.add_out1\[4\] VGND
+ VGND VPWR VPWR _01985_ sky130_fd_sc_hd__nor2b_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07275_ _01926_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09014_ _03498_ _03502_ _02629_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__a21oi_1
XFILLER_132_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09916_ _04188_ _01568_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__or2_1
X_09847_ sha256cu.msg_scheduler.mreg_12\[10\] _04140_ _04146_ _04144_ VGND VGND VPWR
+ VPWR _00425_ sky130_fd_sc_hd__o211a_1
XFILLER_59_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09778_ sha256cu.msg_scheduler.mreg_14\[13\] _04106_ VGND VGND VPWR VPWR _04107_
+ sky130_fd_sc_hd__or2_1
XFILLER_46_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _02081_ _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__xor2_1
XFILLER_73_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _05564_ _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__xor2_1
XFILLER_82_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11671_ _05460_ _05480_ _05479_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__a21boi_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ sha256cu.msg_scheduler.mreg_9\[13\] _04581_ _04591_ _04584_ VGND VGND VPWR
+ VPWR _00761_ sky130_fd_sc_hd__o211a_1
X_14390_ clknet_leaf_15_clk _00904_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13410_ _06706_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10553_ sha256cu.msg_scheduler.mreg_9\[16\] _04548_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__or2_1
X_13341_ _06670_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10484_ sha256cu.msg_scheduler.mreg_8\[19\] _04507_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__or2_1
X_13272_ _06634_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12223_ _06026_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nor2_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12154_ _05747_ _05750_ _05769_ _05962_ _05768_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__a311o_1
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11105_ _04907_ _04961_ _04958_ _04726_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__o211a_2
XFILLER_110_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12085_ _05895_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__nand2_1
XFILLER_77_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11036_ sha256cu.m_pad_pars.block_512\[15\]\[6\] _04781_ _04790_ sha256cu.m_pad_pars.block_512\[11\]\[6\]
+ _04896_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__a221o_1
XFILLER_65_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12987_ sha256cu.m_pad_pars.block_512\[37\]\[2\] _06480_ VGND VGND VPWR VPWR _06483_
+ sky130_fd_sc_hd__and2_1
X_14726_ clknet_leaf_116_clk _01240_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11938_ sha256cu.msg_scheduler.mreg_9\[15\] sha256cu.msg_scheduler.mreg_0\[15\] VGND
+ VGND VPWR VPWR _05756_ sky130_fd_sc_hd__nand2_1
XFILLER_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11869_ _05688_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__nand2_1
XFILLER_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14657_ clknet_leaf_98_clk _01171_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13608_ clknet_leaf_78_clk _00154_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14588_ clknet_leaf_117_clk _01102_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13539_ clknet_leaf_112_clk _00085_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out0\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_13_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07060_ _00457_ _01735_ _01736_ _01741_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__a31o_1
XFILLER_145_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput258 net258 VGND VGND VPWR VPWR cracked sky130_fd_sc_hd__buf_2
XFILLER_99_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07962_ _02574_ _02576_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__xor2_2
X_09701_ sha256cu.iter_processing.w\[12\] _04054_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__or2_1
XFILLER_68_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07893_ _02482_ _02483_ _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__nand3_1
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06913_ _01579_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkinv_2
XFILLER_95_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09632_ _02109_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__buf_4
X_06844_ net19 net22 net21 net25 VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__or4_1
XFILLER_68_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09563_ sha256cu.m_out_digest.f_in\[6\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[6\]
+ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__a22o_1
XFILLER_71_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08514_ _03083_ _03085_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__nand2_1
X_06775_ net257 state\[0\] VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__or2_1
X_09494_ sha256cu.iter_processing.w\[29\] _03089_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__nand2_1
XFILLER_51_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08445_ _02999_ _03001_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__or2b_1
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08376_ _02977_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__xnor2_1
X_07327_ _01969_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07258_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__buf_4
XFILLER_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07189_ _01792_ _01703_ _01598_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__a21o_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13890_ clknet_leaf_24_clk _00436_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12910_ _06441_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__clkbuf_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12841_ sha256cu.m_pad_pars.block_512\[28\]\[6\] _06398_ VGND VGND VPWR VPWR _06405_
+ sky130_fd_sc_hd__and2_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12772_ _06368_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__clkbuf_1
X_11723_ sha256cu.msg_scheduler.mreg_9\[6\] sha256cu.msg_scheduler.mreg_0\[6\] VGND
+ VGND VPWR VPWR _05550_ sky130_fd_sc_hd__or2_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ clknet_leaf_4_clk _01025_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11654_ sha256cu.iter_processing.w\[2\] _05430_ _05484_ _05335_ VGND VGND VPWR VPWR
+ _00900_ sky130_fd_sc_hd__o211a_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ clknet_leaf_9_clk _00956_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10605_ sha256cu.msg_scheduler.mreg_10\[6\] _04574_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__or2_1
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14373_ clknet_leaf_109_clk _00887_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11585_ _04808_ _04912_ _05420_ sha256cu.m_pad_pars.block_512\[48\]\[7\] VGND VGND
+ VPWR VPWR _05421_ sky130_fd_sc_hd__o22a_1
XFILLER_127_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10536_ sha256cu.msg_scheduler.mreg_9\[9\] _04534_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__or2_1
X_13324_ sha256cu.m_pad_pars.block_512\[57\]\[0\] _06660_ VGND VGND VPWR VPWR _06662_
+ sky130_fd_sc_hd__and2_1
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10467_ _04396_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__buf_2
XFILLER_124_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13255_ _06625_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
X_12206_ sha256cu.msg_scheduler.mreg_1\[12\] sha256cu.msg_scheduler.mreg_1\[1\] VGND
+ VGND VPWR VPWR _06013_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10398_ _04396_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__buf_2
XFILLER_89_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13186_ _06588_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12137_ _05916_ _05920_ _05917_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__a21boi_1
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12068_ _05879_ _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__nand2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11019_ sha256cu.data_in_padd\[4\] _01963_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__or2_1
XFILLER_49_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14709_ clknet_leaf_2_clk _01223_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08230_ _02805_ _02797_ _02836_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__and3_1
XANTENNA_390 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08161_ _02739_ _02740_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__and2b_1
XFILLER_146_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08092_ _02684_ _02686_ _02688_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__a21oi_2
X_07112_ _01682_ _01706_ _01787_ _01644_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__a211o_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07043_ _00452_ _01590_ _01583_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__o21ai_2
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08994_ _03482_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__nor2_1
XFILLER_115_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07945_ sha256cu.m_out_digest.b_in\[15\] _02084_ _02559_ VGND VGND VPWR VPWR _02560_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_75_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07876_ _02492_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__inv_2
X_09615_ sha256cu.m_out_digest.g_in\[17\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[17\]
+ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__o22a_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06827_ net68 net71 net70 net73 VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__or4_1
XFILLER_56_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09546_ sha256cu.K\[31\] _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__xnor2_1
X_09477_ _03948_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__nand2_1
X_08428_ _02369_ _03029_ _03030_ _02068_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__a211o_1
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08359_ sha256cu.m_out_digest.e_in\[5\] sha256cu.m_out_digest.e_in\[0\] VGND VGND
+ VPWR VPWR _02963_ sky130_fd_sc_hd__xnor2_2
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11370_ sha256cu.m_pad_pars.block_512\[37\]\[5\] _05165_ _05215_ _05024_ VGND VGND
+ VPWR VPWR _05216_ sky130_fd_sc_hd__a22o_1
XFILLER_20_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10321_ sha256cu.msg_scheduler.mreg_5\[12\] _04407_ _04419_ _04410_ VGND VGND VPWR
+ VPWR _00632_ sky130_fd_sc_hd__o211a_1
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13040_ sha256cu.m_pad_pars.block_512\[40\]\[3\] _06507_ VGND VGND VPWR VPWR _06511_
+ sky130_fd_sc_hd__and2_1
X_10252_ sha256cu.msg_scheduler.mreg_4\[15\] _04367_ _04379_ _04370_ VGND VGND VPWR
+ VPWR _00603_ sky130_fd_sc_hd__o211a_1
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10183_ sha256cu.msg_scheduler.mreg_3\[17\] _04328_ _04340_ _04331_ VGND VGND VPWR
+ VPWR _00573_ sky130_fd_sc_hd__o211a_1
XFILLER_120_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13942_ clknet_leaf_46_clk _00488_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13873_ clknet_leaf_19_clk _00419_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12824_ sha256cu.m_pad_pars.block_512\[27\]\[6\] _06389_ VGND VGND VPWR VPWR _06396_
+ sky130_fd_sc_hd__and2_1
XFILLER_28_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _06359_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11706_ sha256cu.msg_scheduler.mreg_1\[23\] _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__xnor2_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _06322_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11637_ sha256cu.msg_scheduler.mreg_9\[2\] sha256cu.msg_scheduler.mreg_0\[2\] VGND
+ VGND VPWR VPWR _05468_ sky130_fd_sc_hd__nand2_1
X_14425_ clknet_leaf_100_clk _00939_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14356_ clknet_leaf_11_clk _00870_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11568_ _04908_ _05275_ sha256cu.m_pad_pars.block_512\[24\]\[7\] VGND VGND VPWR VPWR
+ _05404_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10519_ sha256cu.msg_scheduler.mreg_8\[1\] _04526_ _04532_ _04530_ VGND VGND VPWR
+ VPWR _00717_ sky130_fd_sc_hd__o211a_1
XFILLER_116_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13307_ sha256cu.m_pad_pars.block_512\[56\]\[0\] _01924_ VGND VGND VPWR VPWR _06653_
+ sky130_fd_sc_hd__and2_1
XFILLER_143_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14287_ clknet_leaf_25_clk _00833_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11499_ sha256cu.m_pad_pars.block_512\[20\]\[2\] _05294_ _05285_ sha256cu.m_pad_pars.block_512\[16\]\[2\]
+ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__a22o_1
X_13238_ _06616_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13169_ _06579_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07730_ _02303_ _02307_ _02350_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__o21a_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07661_ _02281_ _02283_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__xnor2_2
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07592_ _02215_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09400_ _03873_ _03874_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__nand2_1
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09331_ _03777_ _03784_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09262_ _03741_ _03742_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__nor2_1
X_09193_ _03674_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__xnor2_1
X_08213_ sha256cu.iter_processing.w\[22\] _02820_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nor2_1
XFILLER_147_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08144_ _02710_ _02720_ _02753_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__o21ba_1
XFILLER_147_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08075_ _02684_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__xor2_1
XFILLER_115_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07026_ _01593_ _01654_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__nand2_1
XFILLER_121_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08977_ _03466_ _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07928_ sha256cu.K\[13\] _02508_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__a21o_1
XFILLER_68_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07859_ _02470_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__nand2_1
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10870_ sha256cu.m_pad_pars.add_out3\[6\] _01963_ _04738_ _02002_ VGND VGND VPWR
+ VPWR _04740_ sky130_fd_sc_hd__a31o_1
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ _03075_ _03968_ _03967_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12540_ sha256cu.m_pad_pars.block_512\[11\]\[2\] _06241_ VGND VGND VPWR VPWR _06244_
+ sky130_fd_sc_hd__and2_1
X_12471_ _06207_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14210_ clknet_leaf_28_clk _00756_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11422_ _05264_ _04907_ _05265_ sha256cu.m_pad_pars.block_512\[17\]\[7\] VGND VGND
+ VPWR VPWR _05266_ sky130_fd_sc_hd__o22a_1
XFILLER_153_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14141_ clknet_leaf_44_clk _00687_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11353_ sha256cu.data_in_padd\[19\] _04741_ _04742_ _05200_ VGND VGND VPWR VPWR _00882_
+ sky130_fd_sc_hd__a22o_1
X_10304_ _04396_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__buf_2
X_14072_ clknet_leaf_36_clk _00618_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11284_ _04787_ _04993_ _05127_ _05134_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__o211a_2
X_10235_ sha256cu.msg_scheduler.mreg_4\[7\] _04367_ _04369_ _04370_ VGND VGND VPWR
+ VPWR _00595_ sky130_fd_sc_hd__o211a_1
XFILLER_140_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13023_ sha256cu.m_pad_pars.block_512\[39\]\[3\] _06498_ VGND VGND VPWR VPWR _06502_
+ sky130_fd_sc_hd__and2_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10166_ sha256cu.msg_scheduler.mreg_3\[9\] _04328_ _04330_ _04331_ VGND VGND VPWR
+ VPWR _00565_ sky130_fd_sc_hd__o211a_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10097_ sha256cu.msg_scheduler.mreg_3\[12\] _04282_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__or2_1
XFILLER_94_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13925_ clknet_leaf_43_clk _00471_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13856_ clknet_leaf_22_clk _00402_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12807_ sha256cu.m_pad_pars.block_512\[26\]\[6\] _06380_ VGND VGND VPWR VPWR _06387_
+ sky130_fd_sc_hd__and2_1
X_13787_ clknet_leaf_67_clk _00333_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10999_ sha256cu.m_pad_pars.block_512\[31\]\[3\] _04811_ _04861_ _04738_ _04862_
+ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__a221o_1
X_12738_ sha256cu.m_pad_pars.block_512\[22\]\[6\] _06343_ VGND VGND VPWR VPWR _06350_
+ sky130_fd_sc_hd__and2_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _06313_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14408_ clknet_leaf_109_clk _00922_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[24\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14339_ clknet_leaf_111_clk _00853_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out2\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_143_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08900_ _02040_ _03392_ _03393_ _03366_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__o211a_1
XFILLER_112_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09880_ sha256cu.msg_scheduler.mreg_13\[25\] _04160_ VGND VGND VPWR VPWR _04165_
+ sky130_fd_sc_hd__or2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _03325_ _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__xnor2_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08762_ sha256cu.m_out_digest.e_in\[3\] _02732_ _03259_ _03260_ _02258_ VGND VGND
+ VPWR VPWR _00226_ sky130_fd_sc_hd__a221o_1
XFILLER_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07713_ sha256cu.K\[8\] _02319_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__a21boi_1
X_08693_ _03193_ _03194_ sha256cu.K\[0\] VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__a21o_1
X_07644_ _02265_ _02266_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__and2b_1
XFILLER_65_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07575_ sha256cu.m_out_digest.a_in\[27\] _02199_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09314_ _03791_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__or2_1
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09245_ sha256cu.m_out_digest.e_in\[20\] _02439_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__or2_1
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09176_ sha256cu.K\[17\] _03625_ _03624_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__a21o_1
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08127_ sha256cu.iter_processing.w\[19\] _02709_ _02736_ VGND VGND VPWR VPWR _02737_
+ sky130_fd_sc_hd__a21o_1
X_08058_ sha256cu.m_out_digest.b_in\[18\] _02198_ _02669_ VGND VGND VPWR VPWR _02670_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_150_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07009_ _01607_ _01667_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__nor2_2
XFILLER_1_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10020_ _04166_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__buf_2
XFILLER_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput114 hash[201] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xinput103 hash[192] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
Xinput136 hash[221] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput125 hash[211] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xinput147 hash[231] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xinput158 hash[241] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
Xinput169 hash[251] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
X_11971_ _05785_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__nand2_1
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13710_ clknet_leaf_71_clk _00256_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10922_ _04785_ _04786_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__a21o_1
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14690_ clknet_leaf_105_clk _01204_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13641_ clknet_leaf_82_clk _00187_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10853_ _04725_ _01966_ _04723_ _04727_ _01987_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__a32o_1
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10784_ sha256cu.msg_scheduler.mreg_12\[20\] _04679_ VGND VGND VPWR VPWR _04683_
+ sky130_fd_sc_hd__or2_1
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ clknet_leaf_85_clk _00118_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[23\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ sha256cu.m_pad_pars.block_512\[10\]\[2\] _06232_ VGND VGND VPWR VPWR _06235_
+ sky130_fd_sc_hd__and2_1
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12454_ _06198_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__clkbuf_1
X_12385_ sha256cu.m_pad_pars.block_512\[2\]\[1\] _06160_ VGND VGND VPWR VPWR _06162_
+ sky130_fd_sc_hd__and2_1
X_11405_ _04746_ _05248_ sha256cu.m_pad_pars.block_512\[29\]\[7\] VGND VGND VPWR VPWR
+ _05249_ sky130_fd_sc_hd__o21a_1
XFILLER_153_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14124_ clknet_leaf_32_clk _00670_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11336_ sha256cu.m_pad_pars.block_512\[61\]\[2\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[2\]
+ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a22o_1
X_14055_ clknet_leaf_39_clk _00601_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13006_ sha256cu.m_pad_pars.block_512\[38\]\[3\] _06489_ VGND VGND VPWR VPWR _06493_
+ sky130_fd_sc_hd__and2_1
X_11267_ _04933_ _04993_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__o21ai_1
X_10218_ sha256cu.msg_scheduler.mreg_4\[0\] _04354_ _04360_ _04357_ VGND VGND VPWR
+ VPWR _00588_ sky130_fd_sc_hd__o211a_1
X_11198_ sha256cu.m_pad_pars.block_512\[2\]\[4\] _04999_ _05052_ _01921_ VGND VGND
+ VPWR VPWR _05053_ sky130_fd_sc_hd__a22o_1
X_10149_ sha256cu.msg_scheduler.mreg_3\[2\] _04315_ _04321_ _04318_ VGND VGND VPWR
+ VPWR _00558_ sky130_fd_sc_hd__o211a_1
XFILLER_95_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14957_ clknet_leaf_89_clk _01471_ VGND VGND VPWR VPWR sha256cu.K\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_90_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14888_ clknet_leaf_9_clk _01402_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13908_ clknet_leaf_96_clk _00454_ VGND VGND VPWR VPWR sha256cu.counter_iteration\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ clknet_leaf_18_clk _00385_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07360_ sha256cu.m_pad_pars.add_out0\[5\] sha256cu.m_pad_pars.add_out0\[4\] _01992_
+ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__and3_1
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09030_ _03517_ _03518_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__nor2_1
X_07291_ sha256cu.m_pad_pars.add_out0\[3\] sha256cu.m_pad_pars.add_out0\[2\] VGND
+ VGND VPWR VPWR _01935_ sky130_fd_sc_hd__nor2_2
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09932_ _04116_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09863_ sha256cu.msg_scheduler.mreg_12\[17\] _04153_ _04155_ _04144_ VGND VGND VPWR
+ VPWR _00432_ sky130_fd_sc_hd__o211a_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09794_ _01972_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__buf_4
X_08814_ _03309_ _03310_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ sha256cu.K\[3\] _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__xor2_1
XFILLER_100_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ sha256cu.m_out_digest.d_in\[18\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[18\]
+ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__o22a_1
XFILLER_54_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_208 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07627_ sha256cu.K\[5\] _02213_ _02250_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__a21oi_2
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ _02181_ _02182_ _02112_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o21a_1
X_07489_ sha256cu.K\[2\] _02100_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__nand2_1
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09228_ _03708_ _03709_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__nor2_1
XFILLER_148_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09159_ _03620_ _03621_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__nor2_1
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12170_ _05977_ _05978_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__xor2_1
XFILLER_150_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11121_ _04796_ _04824_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__or2_1
XFILLER_1_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11052_ _04704_ _04791_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__or2_4
X_10003_ sha256cu.msg_scheduler.mreg_2\[4\] _04228_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__or2_1
XFILLER_76_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14811_ clknet_leaf_119_clk _01325_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11954_ _05747_ _05750_ _05770_ _05432_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__a31o_1
X_14742_ clknet_leaf_11_clk _01256_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11885_ _05704_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__nand2_1
XFILLER_83_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14673_ clknet_leaf_2_clk _01187_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10905_ _04768_ _04771_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__or2_1
X_13624_ clknet_leaf_63_clk _00170_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10836_ sha256cu.msg_scheduler.counter_iteration\[6\] _04043_ VGND VGND VPWR VPWR
+ _04716_ sky130_fd_sc_hd__nor2_1
X_13555_ clknet_leaf_51_clk _00101_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[6\]
+ sky130_fd_sc_hd__dfxtp_4
X_10767_ sha256cu.msg_scheduler.mreg_11\[12\] _04672_ _04673_ _04662_ VGND VGND VPWR
+ VPWR _00824_ sky130_fd_sc_hd__o211a_1
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10698_ sha256cu.msg_scheduler.mreg_10\[14\] _04633_ _04634_ _04623_ VGND VGND VPWR
+ VPWR _00794_ sky130_fd_sc_hd__o211a_1
XFILLER_12_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12506_ sha256cu.m_pad_pars.block_512\[9\]\[2\] _06223_ VGND VGND VPWR VPWR _06226_
+ sky130_fd_sc_hd__and2_1
X_13486_ _06755_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_1
X_12437_ _06189_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14107_ clknet_leaf_36_clk _00653_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12368_ _06153_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12299_ _06080_ _06082_ _06079_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__a21boi_1
X_11319_ sha256cu.m_pad_pars.block_512\[45\]\[0\] _05126_ _05133_ _05169_ VGND VGND
+ VPWR VPWR _05170_ sky130_fd_sc_hd__a211o_1
XFILLER_4_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14038_ clknet_leaf_39_clk _00584_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06860_ _01554_ _01555_ _01556_ _01557_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__or4_2
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06791_ net182 net185 net184 net187 VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__or4_1
XFILLER_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08530_ _03123_ _03128_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__nor2_1
XFILLER_48_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08461_ _03060_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07412_ _02019_ _02020_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__and2b_1
XFILLER_51_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08392_ _02994_ _02995_ _02161_ _02070_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__a2bb2o_1
X_07343_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__buf_4
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07274_ sha256cu.m_pad_pars.block_512\[63\]\[1\] _01924_ VGND VGND VPWR VPWR _01926_
+ sky130_fd_sc_hd__and2_1
XFILLER_148_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09013_ _03498_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__or2_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09915_ sha256cu.counter_iteration\[6\] VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__buf_2
X_09846_ sha256cu.msg_scheduler.mreg_13\[10\] _04134_ VGND VGND VPWR VPWR _04146_
+ sky130_fd_sc_hd__or2_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _04053_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__clkbuf_2
XFILLER_74_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06989_ _01617_ _01661_ _01673_ _01676_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__a31o_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _03226_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nand2_1
XFILLER_100_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ sha256cu.m_out_digest.d_in\[5\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[5\]
+ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__o22a_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11670_ _05497_ _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__xnor2_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10621_ sha256cu.msg_scheduler.mreg_10\[13\] _04588_ VGND VGND VPWR VPWR _04591_
+ sky130_fd_sc_hd__or2_1
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10552_ sha256cu.msg_scheduler.mreg_8\[15\] _04540_ _04551_ _04543_ VGND VGND VPWR
+ VPWR _00731_ sky130_fd_sc_hd__o211a_1
X_13340_ sha256cu.m_pad_pars.block_512\[58\]\[0\] _06660_ VGND VGND VPWR VPWR _06670_
+ sky130_fd_sc_hd__and2_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13271_ sha256cu.m_pad_pars.block_512\[53\]\[7\] _05235_ _01965_ VGND VGND VPWR VPWR
+ _06634_ sky130_fd_sc_hd__mux2_1
X_10483_ sha256cu.msg_scheduler.mreg_7\[18\] _04500_ _04511_ _04503_ VGND VGND VPWR
+ VPWR _00702_ sky130_fd_sc_hd__o211a_1
X_12222_ _05967_ _06027_ _06028_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__o21a_1
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12153_ _05886_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__or2_1
XFILLER_151_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12084_ sha256cu.msg_scheduler.mreg_9\[21\] sha256cu.msg_scheduler.mreg_0\[21\] VGND
+ VGND VPWR VPWR _05896_ sky130_fd_sc_hd__nand2_1
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11104_ _04959_ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__nor2_4
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11035_ sha256cu.m_pad_pars.block_512\[59\]\[6\] _04829_ _04833_ sha256cu.m_pad_pars.block_512\[55\]\[6\]
+ _04895_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__a221o_1
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12986_ _06482_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14725_ clknet_leaf_100_clk _01239_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11937_ sha256cu.msg_scheduler.mreg_9\[15\] sha256cu.msg_scheduler.mreg_0\[15\] VGND
+ VGND VPWR VPWR _05755_ sky130_fd_sc_hd__or2_1
XFILLER_45_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11868_ sha256cu.msg_scheduler.mreg_9\[12\] sha256cu.msg_scheduler.mreg_0\[12\] VGND
+ VGND VPWR VPWR _05689_ sky130_fd_sc_hd__nand2_1
X_14656_ clknet_leaf_96_clk _01170_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11799_ _05621_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__nand2_1
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13607_ clknet_leaf_79_clk _00153_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14587_ clknet_leaf_118_clk _01101_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10819_ _04702_ _04705_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__nor2_1
X_13538_ clknet_leaf_109_clk _00035_ VGND VGND VPWR VPWR state\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13469_ _06730_ _06744_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__and2_1
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput259 net259 VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_2
XFILLER_114_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07961_ _02523_ _02533_ _02575_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__o21bai_2
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09700_ sha256cu.msg_scheduler.mreg_14\[11\] _04060_ _04062_ _04050_ VGND VGND VPWR
+ VPWR _00362_ sky130_fd_sc_hd__o211a_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06912_ _01601_ _01603_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__nor2_2
X_07892_ sha256cu.K\[13\] _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06843_ net15 net18 net17 net20 VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__or4_2
XFILLER_95_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09631_ sha256cu.m_out_digest.g_in\[31\] _04037_ _04036_ sha256cu.m_out_digest.f_in\[31\]
+ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__a22o_1
X_09562_ sha256cu.m_out_digest.f_in\[5\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[5\]
+ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__a22o_1
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08513_ _03097_ _03099_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__nor2_1
X_09493_ sha256cu.iter_processing.w\[29\] _03089_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__or2_1
XFILLER_24_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08444_ _03043_ _03045_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08375_ sha256cu.iter_processing.w\[25\] _02940_ _02978_ VGND VGND VPWR VPWR _02979_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_11_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07326_ _01938_ _01960_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__or2_2
XFILLER_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07257_ _01564_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__clkinv_4
XFILLER_133_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07188_ _01808_ _01650_ _01627_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__or3b_1
XFILLER_132_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09829_ sha256cu.msg_scheduler.mreg_12\[2\] _04126_ _04136_ _04130_ VGND VGND VPWR
+ VPWR _00417_ sky130_fd_sc_hd__o211a_1
XFILLER_86_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12840_ _06404_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__clkbuf_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12771_ sha256cu.m_pad_pars.block_512\[24\]\[5\] _06362_ VGND VGND VPWR VPWR _06368_
+ sky130_fd_sc_hd__and2_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ sha256cu.iter_processing.w\[5\] _05430_ _05549_ _05335_ VGND VGND VPWR VPWR
+ _00903_ sky130_fd_sc_hd__o211a_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ clknet_leaf_109_clk _01024_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11653_ sha256cu.data_in_padd\[2\] _05448_ _05483_ _05463_ VGND VGND VPWR VPWR _05484_
+ sky130_fd_sc_hd__a211o_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ clknet_leaf_11_clk _00955_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10604_ _04580_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__clkbuf_4
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14372_ clknet_leaf_110_clk _00886_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_13323_ _06661_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__clkbuf_1
X_11584_ _04824_ _05136_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__nor2_1
X_10535_ sha256cu.msg_scheduler.mreg_8\[8\] _04540_ _04541_ _04530_ VGND VGND VPWR
+ VPWR _00724_ sky130_fd_sc_hd__o211a_1
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10466_ sha256cu.msg_scheduler.mreg_8\[11\] _04494_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__or2_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13254_ sha256cu.m_pad_pars.block_512\[52\]\[7\] _05415_ _06542_ VGND VGND VPWR VPWR
+ _06625_ sky130_fd_sc_hd__mux2_1
X_12205_ _06010_ _06011_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__nand2_1
XFILLER_6_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13185_ sha256cu.m_pad_pars.block_512\[48\]\[7\] _05421_ _06542_ VGND VGND VPWR VPWR
+ _06588_ sky130_fd_sc_hd__mux2_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10397_ sha256cu.msg_scheduler.mreg_7\[13\] _04455_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__or2_1
XFILLER_123_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12136_ _05943_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__xor2_1
XFILLER_69_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12067_ _05876_ _05878_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__or2_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11018_ _04876_ _04878_ _04879_ _04880_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__or4_2
XFILLER_65_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12969_ _06473_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__clkbuf_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14708_ clknet_leaf_5_clk _01222_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_380 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14639_ clknet_leaf_9_clk _01153_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_391 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08160_ _02768_ _02769_ _02273_ _02070_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_118_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07111_ _01649_ _01696_ _01603_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__o21a_1
X_08091_ sha256cu.K\[18\] _02691_ _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__a21boi_2
XFILLER_146_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07042_ _01617_ _01720_ _01724_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__a21o_1
XFILLER_130_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08993_ sha256cu.iter_processing.w\[12\] _02446_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__and2_1
XFILLER_130_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07944_ sha256cu.m_out_digest.b_in\[15\] _02084_ sha256cu.m_out_digest.c_in\[15\]
+ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__a21o_1
X_07875_ sha256cu.m_out_digest.e_in\[24\] _02491_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__xnor2_4
XFILLER_56_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06826_ net59 net62 net61 net64 VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__or4_2
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09614_ sha256cu.m_out_digest.g_in\[16\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[16\]
+ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__o22a_1
XFILLER_83_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09545_ _03119_ _03987_ _03986_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__a21oi_1
X_09476_ _03916_ _03917_ _03949_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08427_ sha256cu.m_out_digest.a_in\[27\] _02629_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__and2_1
XFILLER_12_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08358_ sha256cu.m_out_digest.h_in\[26\] _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__xnor2_1
X_08289_ sha256cu.m_out_digest.e_in\[30\] _02894_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__xnor2_4
X_07309_ sha256cu.m_pad_pars.add_512_block\[3\] sha256cu.m_pad_pars.add_512_block\[2\]
+ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__nand2b_2
XFILLER_20_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10320_ sha256cu.msg_scheduler.mreg_6\[12\] _04415_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__or2_1
XFILLER_106_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10251_ sha256cu.msg_scheduler.mreg_5\[15\] _04374_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__or2_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10182_ sha256cu.msg_scheduler.mreg_4\[17\] _04335_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__or2_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13941_ clknet_leaf_46_clk _00487_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13872_ clknet_leaf_18_clk _00418_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12823_ _06395_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ sha256cu.m_pad_pars.block_512\[23\]\[5\] _06353_ VGND VGND VPWR VPWR _06359_
+ sky130_fd_sc_hd__and2_1
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11705_ sha256cu.msg_scheduler.mreg_1\[12\] sha256cu.msg_scheduler.mreg_1\[8\] VGND
+ VGND VPWR VPWR _05533_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ sha256cu.m_pad_pars.block_512\[19\]\[5\] _06316_ VGND VGND VPWR VPWR _06322_
+ sky130_fd_sc_hd__and2_1
XFILLER_15_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11636_ _05456_ _05458_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__nand2_1
X_14424_ clknet_leaf_117_clk _00938_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14355_ clknet_leaf_14_clk _00869_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11567_ _05278_ _05297_ _05400_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__a31o_1
X_10518_ sha256cu.msg_scheduler.mreg_9\[1\] _04520_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__or2_1
X_14286_ clknet_leaf_24_clk _00832_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13306_ _06652_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13237_ sha256cu.m_pad_pars.block_512\[51\]\[7\] _04932_ _06542_ VGND VGND VPWR VPWR
+ _06616_ sky130_fd_sc_hd__mux2_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11498_ sha256cu.m_pad_pars.block_512\[12\]\[2\] _05299_ _05304_ sha256cu.m_pad_pars.block_512\[36\]\[2\]
+ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__a221o_1
X_10449_ sha256cu.msg_scheduler.mreg_7\[3\] _04487_ _04492_ _04490_ VGND VGND VPWR
+ VPWR _00687_ sky130_fd_sc_hd__o211a_1
XFILLER_112_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13168_ sha256cu.m_pad_pars.block_512\[47\]\[7\] _04919_ _06542_ VGND VGND VPWR VPWR
+ _06579_ sky130_fd_sc_hd__mux2_1
X_12119_ _05904_ _05906_ _05902_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__a21oi_1
X_13099_ _01964_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__buf_4
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07660_ _02228_ _02240_ _02282_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__o21ba_1
X_07591_ _02178_ _02180_ _02183_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__o21a_1
X_09330_ _03807_ _03808_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__nor2_1
XFILLER_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09261_ _03736_ _03740_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__and2_1
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08212_ _02818_ _02819_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__xnor2_1
X_09192_ _02675_ _03644_ _03645_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__a21boi_1
XFILLER_135_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08143_ _02717_ _02719_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__nor2_1
XFILLER_147_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08074_ _02641_ _02651_ _02685_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__o21bai_2
XFILLER_134_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07025_ _01709_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08976_ _03431_ _03434_ _03433_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07927_ _02505_ _02507_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__nor2_1
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07858_ _02329_ _02472_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__o21ba_1
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07789_ _02394_ _02396_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__or2b_1
XFILLER_84_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06809_ net135 net138 net137 net140 VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__or4_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09528_ _03998_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__nor2_1
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09459_ _03001_ _03900_ _03899_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__a21boi_1
X_12470_ sha256cu.m_pad_pars.block_512\[7\]\[1\] _06205_ VGND VGND VPWR VPWR _06207_
+ sky130_fd_sc_hd__and2_1
XFILLER_40_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11421_ _04807_ _05004_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__nor2_1
XFILLER_126_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14140_ clknet_leaf_36_clk _00686_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11352_ _05192_ _05194_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__or3_1
XFILLER_153_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10303_ sha256cu.msg_scheduler.mreg_6\[5\] _04401_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__or2_1
XFILLER_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14071_ clknet_leaf_36_clk _00617_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11283_ sha256cu.m_pad_pars.add_out1\[3\] sha256cu.m_pad_pars.add_out1\[2\] VGND
+ VGND VPWR VPWR _05134_ sky130_fd_sc_hd__nor2_2
X_10234_ _04263_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__buf_2
XFILLER_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13022_ _06501_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__clkbuf_1
X_10165_ _04263_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__buf_2
XFILLER_105_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10096_ sha256cu.msg_scheduler.mreg_2\[11\] _04288_ _04290_ _04291_ VGND VGND VPWR
+ VPWR _00535_ sky130_fd_sc_hd__o211a_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13924_ clknet_leaf_44_clk _00470_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ clknet_leaf_22_clk _00401_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12806_ _06386_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13786_ clknet_leaf_67_clk _00332_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10998_ sha256cu.m_pad_pars.block_512\[59\]\[3\] _04829_ _04833_ sha256cu.m_pad_pars.block_512\[55\]\[3\]
+ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__a22o_1
X_12737_ _06349_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__clkbuf_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12668_ sha256cu.m_pad_pars.block_512\[18\]\[5\] _06307_ VGND VGND VPWR VPWR _06313_
+ sky130_fd_sc_hd__and2_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11619_ _05449_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nand2_1
X_14407_ clknet_leaf_77_clk _00921_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[23\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12599_ _06276_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14338_ clknet_leaf_105_clk _00852_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.counter_iteration\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14269_ clknet_leaf_18_clk _00815_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _02196_ _03293_ _03292_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08761_ _03237_ _03258_ _02515_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__o21a_1
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07712_ _02316_ _02318_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__or2b_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08692_ sha256cu.iter_processing.w\[0\] _02020_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__or2_1
X_07643_ _02262_ _02263_ _02264_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a21o_1
XFILLER_81_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07574_ _02198_ sha256cu.m_out_digest.a_in\[7\] VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__xnor2_1
X_09313_ _03789_ _03790_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__and2_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_60_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
X_09244_ _03719_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__xnor2_1
X_09175_ _03657_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__and2_1
XFILLER_147_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08126_ _02707_ _02708_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__and2b_1
XFILLER_134_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08057_ sha256cu.m_out_digest.b_in\[18\] _02198_ sha256cu.m_out_digest.c_in\[18\]
+ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07008_ _01679_ _01683_ _01686_ _01693_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__a31o_1
XFILLER_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput104 hash[193] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_2
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput115 hash[202] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
Xinput126 hash[212] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
X_08959_ _03437_ _03436_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__or2b_1
XFILLER_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput148 hash[232] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xinput137 hash[222] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xinput159 hash[242] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
X_11970_ sha256cu.msg_scheduler.mreg_14\[26\] _05786_ VGND VGND VPWR VPWR _05787_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_91_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10921_ _04751_ _04787_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__nor2_1
XFILLER_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13640_ clknet_leaf_78_clk _00186_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10852_ sha256cu.m_pad_pars.add_out2\[3\] sha256cu.m_pad_pars.add_out2\[2\] _04726_
+ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__and3_1
X_10783_ sha256cu.msg_scheduler.mreg_11\[19\] _04672_ _04682_ _04675_ VGND VGND VPWR
+ VPWR _00831_ sky130_fd_sc_hd__o211a_1
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ clknet_leaf_86_clk _00117_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _06234_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12453_ sha256cu.m_pad_pars.block_512\[6\]\[1\] _06196_ VGND VGND VPWR VPWR _06198_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12384_ _06161_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_1
X_11404_ _01941_ _04776_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__or2_2
XFILLER_153_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14123_ clknet_leaf_32_clk _00669_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11335_ sha256cu.m_pad_pars.block_512\[17\]\[2\] _05138_ _05158_ sha256cu.m_pad_pars.block_512\[21\]\[2\]
+ _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__a221o_1
XFILLER_153_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14054_ clknet_leaf_40_clk _00600_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11266_ _01944_ _04699_ _05117_ sha256cu.m_pad_pars.block_512\[2\]\[7\] VGND VGND
+ VPWR VPWR _05118_ sky130_fd_sc_hd__a31o_1
XFILLER_141_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10217_ sha256cu.msg_scheduler.mreg_5\[0\] _04348_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__or2_1
XFILLER_106_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13005_ _06492_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11197_ sha256cu.m_pad_pars.block_512\[62\]\[4\] _04984_ _04982_ sha256cu.m_pad_pars.block_512\[58\]\[4\]
+ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__a22o_1
X_10148_ sha256cu.msg_scheduler.mreg_4\[2\] _04308_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__or2_1
XFILLER_94_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10079_ _01566_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14956_ clknet_leaf_89_clk _01470_ VGND VGND VPWR VPWR sha256cu.K\[29\] sky130_fd_sc_hd__dfxtp_1
X_13907_ clknet_leaf_97_clk _00453_ VGND VGND VPWR VPWR sha256cu.counter_iteration\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14887_ clknet_leaf_123_clk _01401_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13838_ clknet_leaf_17_clk _00384_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13769_ clknet_leaf_82_clk _00315_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_42_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07290_ _01934_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09931_ sha256cu.msg_scheduler.mreg_1\[5\] _04174_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__or2_1
XFILLER_116_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09862_ sha256cu.msg_scheduler.mreg_13\[17\] _04147_ VGND VGND VPWR VPWR _04155_
+ sky130_fd_sc_hd__or2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08813_ _03282_ _03284_ _03286_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__o21ba_1
XFILLER_85_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09793_ sha256cu.msg_scheduler.mreg_14\[20\] _04106_ VGND VGND VPWR VPWR _04115_
+ sky130_fd_sc_hd__or2_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _03241_ _03242_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__nand2_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ sha256cu.m_out_digest.d_in\[17\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[17\]
+ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__o22a_1
XFILLER_54_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_209 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07626_ _02210_ _02212_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__nor2_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07557_ _02181_ _02182_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_33_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_139_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07488_ _02096_ _02099_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__or2_1
XFILLER_42_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09227_ _03703_ _03707_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__and2_1
XFILLER_10_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09158_ _03632_ _03633_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__nand2_1
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09089_ _03574_ _03575_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__xnor2_1
X_08109_ _02717_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11120_ _01952_ _04969_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__or2_1
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11051_ _04907_ _04779_ _04910_ sha256cu.m_pad_pars.block_512\[31\]\[7\] VGND VGND
+ VPWR VPWR _04911_ sky130_fd_sc_hd__o22a_1
X_10002_ sha256cu.msg_scheduler.mreg_1\[3\] _04234_ _04236_ _04237_ VGND VGND VPWR
+ VPWR _00495_ sky130_fd_sc_hd__o211a_1
XFILLER_130_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14810_ clknet_leaf_118_clk _01324_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11953_ _05747_ _05750_ _05770_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14741_ clknet_leaf_3_clk _01255_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11884_ _05702_ _05703_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__nand2_1
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10904_ _01953_ _04752_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__or2_2
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14672_ clknet_leaf_2_clk _01186_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13623_ clknet_leaf_63_clk _00169_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10835_ sha256cu.msg_scheduler.temp_case _04190_ sha256cu.msg_scheduler.counter_iteration\[0\]
+ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_24_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
X_13554_ clknet_leaf_51_clk _00100_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[5\]
+ sky130_fd_sc_hd__dfxtp_4
X_10766_ sha256cu.msg_scheduler.mreg_12\[12\] _04666_ VGND VGND VPWR VPWR _04673_
+ sky130_fd_sc_hd__or2_1
X_10697_ sha256cu.msg_scheduler.mreg_11\[14\] _04627_ VGND VGND VPWR VPWR _04634_
+ sky130_fd_sc_hd__or2_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13485_ _06730_ _06754_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__and2_1
X_12505_ _06225_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12436_ sha256cu.m_pad_pars.block_512\[5\]\[1\] _06187_ VGND VGND VPWR VPWR _06189_
+ sky130_fd_sc_hd__and2_1
X_14106_ clknet_leaf_36_clk _00652_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12367_ sha256cu.m_pad_pars.block_512\[1\]\[0\] _06152_ VGND VGND VPWR VPWR _06153_
+ sky130_fd_sc_hd__and2_1
X_12298_ _06099_ _06100_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__xor2_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11318_ _05143_ _05148_ _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__or3_1
X_14037_ clknet_leaf_39_clk _00583_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11249_ _04908_ _04973_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__nand2_1
XFILLER_68_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06790_ net167 net176 net175 net178 VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__or4_1
X_14939_ clknet_leaf_91_clk _01453_ VGND VGND VPWR VPWR sha256cu.K\[12\] sky130_fd_sc_hd__dfxtp_4
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08460_ sha256cu.iter_processing.w\[27\] _03009_ _03061_ VGND VGND VPWR VPWR _03062_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_36_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07411_ _02037_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__buf_4
X_08391_ _02988_ _02993_ _02478_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__a21o_1
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
X_07342_ _01964_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__buf_4
XFILLER_16_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07273_ _01925_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09012_ _03391_ _03444_ _03499_ _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__o31a_2
XFILLER_117_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09914_ _04187_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09845_ sha256cu.msg_scheduler.mreg_12\[9\] _04140_ _04145_ _04144_ VGND VGND VPWR
+ VPWR _00424_ sky130_fd_sc_hd__o211a_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09776_ sha256cu.msg_scheduler.mreg_13\[12\] _04099_ _04105_ _04103_ VGND VGND VPWR
+ VPWR _00395_ sky130_fd_sc_hd__o211a_1
X_06988_ _01674_ _01675_ _01596_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__o21a_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ sha256cu.m_out_digest.h_in\[2\] sha256cu.m_out_digest.d_in\[2\] VGND VGND
+ VPWR VPWR _03227_ sky130_fd_sc_hd__or2_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ sha256cu.m_out_digest.d_in\[4\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[4\]
+ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__o22a_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ sha256cu.m_out_digest.a_in\[19\] VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08589_ sha256cu.m_out_digest.b_in\[11\] _02370_ _02110_ sha256cu.m_out_digest.a_in\[11\]
+ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__o22a_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10620_ sha256cu.msg_scheduler.mreg_9\[12\] _04581_ _04590_ _04584_ VGND VGND VPWR
+ VPWR _00760_ sky130_fd_sc_hd__o211a_1
X_10551_ sha256cu.msg_scheduler.mreg_9\[15\] _04548_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__or2_1
X_10482_ sha256cu.msg_scheduler.mreg_8\[18\] _04507_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__or2_1
X_13270_ _06633_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
X_12221_ _05981_ _06004_ _06003_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__a21o_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12152_ _05934_ _05935_ _05956_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__nand3_1
XFILLER_151_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12083_ sha256cu.msg_scheduler.mreg_9\[21\] sha256cu.msg_scheduler.mreg_0\[21\] VGND
+ VGND VPWR VPWR _05895_ sky130_fd_sc_hd__or2_1
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11103_ _04769_ _04961_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__nor2_1
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11034_ sha256cu.m_pad_pars.block_512\[35\]\[6\] _04818_ _04894_ _04738_ VGND VGND
+ VPWR VPWR _04895_ sky130_fd_sc_hd__a22o_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12985_ sha256cu.m_pad_pars.block_512\[37\]\[1\] _06480_ VGND VGND VPWR VPWR _06482_
+ sky130_fd_sc_hd__and2_1
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11936_ sha256cu.iter_processing.w\[14\] _05666_ _05754_ _05640_ VGND VGND VPWR VPWR
+ _00912_ sky130_fd_sc_hd__o211a_1
X_14724_ clknet_leaf_100_clk _01238_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11867_ sha256cu.msg_scheduler.mreg_9\[12\] sha256cu.msg_scheduler.mreg_0\[12\] VGND
+ VGND VPWR VPWR _05688_ sky130_fd_sc_hd__or2_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14655_ clknet_leaf_98_clk _01169_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11798_ sha256cu.msg_scheduler.mreg_9\[9\] sha256cu.msg_scheduler.mreg_0\[9\] VGND
+ VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nand2_1
X_13606_ clknet_leaf_80_clk _00152_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14586_ clknet_leaf_118_clk _01100_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10818_ _04704_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__clkbuf_4
X_10749_ sha256cu.msg_scheduler.mreg_11\[4\] _04659_ _04663_ _04662_ VGND VGND VPWR
+ VPWR _00816_ sky130_fd_sc_hd__o211a_1
X_13537_ clknet_leaf_109_clk _00034_ VGND VGND VPWR VPWR state\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13468_ sha256cu.K\[14\] _06714_ _06719_ _00041_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__a22o_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12419_ sha256cu.m_pad_pars.block_512\[4\]\[1\] _06178_ VGND VGND VPWR VPWR _06180_
+ sky130_fd_sc_hd__and2_1
X_13399_ sha256cu.m_pad_pars.block_512\[61\]\[4\] _06693_ VGND VGND VPWR VPWR _06701_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07960_ _02530_ _02532_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__nor2_1
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_06911_ _01602_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_4
X_07891_ _02505_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__xor2_1
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06842_ net6 net9 net8 net11 VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__or4_1
X_09630_ sha256cu.m_out_digest.g_in\[30\] _04037_ _04036_ sha256cu.m_out_digest.f_in\[30\]
+ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__a22o_1
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09561_ sha256cu.m_out_digest.f_in\[4\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[4\]
+ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__a22o_1
XFILLER_67_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08512_ _03075_ _03103_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nor2_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09492_ _03963_ _03964_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__or2_1
XFILLER_24_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08443_ sha256cu.m_out_digest.e_in\[21\] _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__xnor2_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08374_ _02938_ _02939_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__and2b_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07325_ sha256cu.m_pad_pars.add_out1\[3\] sha256cu.m_pad_pars.add_out1\[2\] VGND
+ VGND VPWR VPWR _01968_ sky130_fd_sc_hd__nand2_1
XFILLER_32_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07256_ state\[2\] VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__inv_2
XFILLER_137_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07187_ _01679_ _01848_ _01850_ _01853_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__a31o_1
XFILLER_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09828_ sha256cu.msg_scheduler.mreg_13\[2\] _04134_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__or2_1
XFILLER_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09759_ sha256cu.msg_scheduler.mreg_14\[5\] _04093_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__or2_1
XFILLER_46_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _06367_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__clkbuf_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ sha256cu.data_in_padd\[5\] _05448_ _05548_ _05463_ VGND VGND VPWR VPWR _05549_
+ sky130_fd_sc_hd__a211o_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11652_ _05465_ _05481_ _05482_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__nor3_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ clknet_leaf_9_clk _00954_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10603_ _04043_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__clkbuf_4
X_14371_ clknet_leaf_77_clk _00885_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13322_ sha256cu.m_pad_pars.block_512\[56\]\[7\] _06660_ VGND VGND VPWR VPWR _06661_
+ sky130_fd_sc_hd__and2_1
X_11583_ sha256cu.m_pad_pars.block_512\[60\]\[7\] _01997_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[7\]
+ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__a22o_1
X_10534_ sha256cu.msg_scheduler.mreg_9\[8\] _04534_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__or2_1
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10465_ sha256cu.msg_scheduler.mreg_7\[10\] _04500_ _04501_ _04490_ VGND VGND VPWR
+ VPWR _00694_ sky130_fd_sc_hd__o211a_1
XFILLER_109_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13253_ _06624_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
X_10396_ sha256cu.msg_scheduler.mreg_6\[12\] _04461_ _04462_ _04451_ VGND VGND VPWR
+ VPWR _00664_ sky130_fd_sc_hd__o211a_1
X_12204_ sha256cu.msg_scheduler.mreg_9\[26\] sha256cu.msg_scheduler.mreg_0\[26\] VGND
+ VGND VPWR VPWR _06011_ sky130_fd_sc_hd__nand2_1
X_13184_ _06587_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12135_ sha256cu.msg_scheduler.mreg_1\[30\] _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12066_ _05876_ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__nand2_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11017_ sha256cu.m_pad_pars.block_512\[15\]\[4\] _04781_ _04800_ sha256cu.m_pad_pars.block_512\[39\]\[4\]
+ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__a22o_1
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12968_ sha256cu.m_pad_pars.block_512\[36\]\[1\] _06471_ VGND VGND VPWR VPWR _06473_
+ sky130_fd_sc_hd__and2_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11919_ _05736_ _05737_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__or2_1
XANTENNA_370 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14707_ clknet_leaf_5_clk _01221_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12899_ sha256cu.m_pad_pars.block_512\[32\]\[1\] _06434_ VGND VGND VPWR VPWR _06436_
+ sky130_fd_sc_hd__and2_1
XANTENNA_381 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14638_ clknet_leaf_108_clk _01152_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_392 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14569_ clknet_leaf_16_clk _01083_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_07110_ _01679_ _01782_ _01786_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__a21o_1
XFILLER_118_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08090_ _02690_ _02666_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__or2b_1
X_07041_ _01722_ _01723_ _01584_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__a21oi_1
XFILLER_133_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08992_ sha256cu.iter_processing.w\[12\] _02446_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__nor2_1
XFILLER_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07943_ sha256cu.iter_processing.w\[14\] _02522_ _02557_ VGND VGND VPWR VPWR _02558_
+ sky130_fd_sc_hd__a21o_1
X_07874_ sha256cu.m_out_digest.e_in\[19\] sha256cu.m_out_digest.e_in\[6\] VGND VGND
+ VPWR VPWR _02491_ sky130_fd_sc_hd__xnor2_2
X_09613_ sha256cu.m_out_digest.g_in\[15\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[15\]
+ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__o22a_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06825_ net63 net66 net65 net69 VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__or4_4
XFILLER_141_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09544_ _03157_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__xor2_1
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09475_ _03915_ _03914_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__or2b_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08426_ _03026_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__xor2_1
XFILLER_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08357_ _02232_ _02960_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08288_ sha256cu.m_out_digest.e_in\[17\] sha256cu.m_out_digest.e_in\[3\] VGND VGND
+ VPWR VPWR _02894_ sky130_fd_sc_hd__xnor2_2
X_07308_ _01951_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07239_ _01724_ _01897_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__or2_1
X_10250_ sha256cu.msg_scheduler.mreg_4\[14\] _04367_ _04378_ _04370_ VGND VGND VPWR
+ VPWR _00602_ sky130_fd_sc_hd__o211a_1
XFILLER_133_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10181_ sha256cu.msg_scheduler.mreg_3\[16\] _04328_ _04339_ _04331_ VGND VGND VPWR
+ VPWR _00572_ sky130_fd_sc_hd__o211a_1
XFILLER_105_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13940_ clknet_leaf_49_clk _00486_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13871_ clknet_leaf_21_clk _00417_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12822_ sha256cu.m_pad_pars.block_512\[27\]\[5\] _06389_ VGND VGND VPWR VPWR _06395_
+ sky130_fd_sc_hd__and2_1
XFILLER_27_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _06358_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11704_ _05530_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__nand2_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _06321_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14423_ clknet_leaf_120_clk _00937_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11635_ _05454_ _05455_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__or2_1
X_14354_ clknet_leaf_14_clk _00868_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11566_ _05293_ _05297_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and3_1
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10517_ sha256cu.msg_scheduler.mreg_8\[0\] _04526_ _04531_ _04530_ VGND VGND VPWR
+ VPWR _00716_ sky130_fd_sc_hd__o211a_1
X_14285_ clknet_leaf_24_clk _00831_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13305_ sha256cu.m_pad_pars.block_512\[55\]\[7\] _06644_ VGND VGND VPWR VPWR _06652_
+ sky130_fd_sc_hd__and2_1
X_13236_ _06615_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_1
X_11497_ sha256cu.m_pad_pars.block_512\[4\]\[2\] _05313_ _05320_ sha256cu.m_pad_pars.block_512\[40\]\[2\]
+ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__a22o_1
XFILLER_6_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10448_ sha256cu.msg_scheduler.mreg_8\[3\] _04481_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__or2_1
X_10379_ sha256cu.msg_scheduler.mreg_7\[5\] _04441_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__or2_1
XFILLER_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13167_ _06578_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__clkbuf_1
X_12118_ _05927_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__nand2_1
XFILLER_69_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13098_ _06541_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12049_ _05838_ _05841_ _05861_ _05465_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__a31o_1
XFILLER_1_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07590_ _02186_ _02214_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__xor2_1
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09260_ _03736_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__nor2_1
X_08211_ sha256cu.m_out_digest.g_in\[22\] sha256cu.m_out_digest.f_in\[22\] sha256cu.m_out_digest.e_in\[22\]
+ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__mux2_2
XFILLER_61_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09191_ _02712_ _03673_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__xor2_1
X_08142_ _02742_ _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__xor2_2
XFILLER_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08073_ _02648_ _02650_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__nor2_1
X_07024_ _01699_ _01708_ _01570_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__mux2_1
XFILLER_103_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08975_ _03464_ _03465_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07926_ sha256cu.K\[14\] _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__xnor2_2
XFILLER_111_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07857_ _02436_ _02473_ _02471_ _02405_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__a221o_1
XFILLER_72_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07788_ sha256cu.m_out_digest.a_in\[10\] _02370_ _02110_ _02407_ VGND VGND VPWR VPWR
+ _00105_ sky130_fd_sc_hd__o22a_1
XFILLER_84_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06808_ net170 net173 net172 _01505_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__or4_2
X_09527_ _03963_ _03970_ _03997_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__nor3_1
XFILLER_71_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09458_ _03045_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__xor2_1
XFILLER_24_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09389_ _03832_ _03840_ _03865_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__and3_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08409_ _03005_ _03010_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__or2_1
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11420_ _01940_ _01941_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__or2_1
XFILLER_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11351_ sha256cu.m_pad_pars.block_512\[45\]\[3\] _05126_ _05132_ sha256cu.m_pad_pars.block_512\[41\]\[3\]
+ _05198_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__a221o_1
XFILLER_137_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10302_ sha256cu.msg_scheduler.mreg_5\[4\] _04407_ _04408_ _04397_ VGND VGND VPWR
+ VPWR _00624_ sky130_fd_sc_hd__o211a_1
XFILLER_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14070_ clknet_leaf_38_clk _00616_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11282_ sha256cu.m_pad_pars.block_512\[13\]\[0\] _05128_ _05132_ sha256cu.m_pad_pars.block_512\[41\]\[0\]
+ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__a22o_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10233_ sha256cu.msg_scheduler.mreg_5\[7\] _04361_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__or2_1
XFILLER_105_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13021_ sha256cu.m_pad_pars.block_512\[39\]\[2\] _06498_ VGND VGND VPWR VPWR _06501_
+ sky130_fd_sc_hd__and2_1
X_10164_ sha256cu.msg_scheduler.mreg_4\[9\] _04322_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__or2_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10095_ _04263_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__buf_2
XFILLER_120_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13923_ clknet_leaf_44_clk _00469_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13854_ clknet_leaf_17_clk _00400_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12805_ sha256cu.m_pad_pars.block_512\[26\]\[5\] _06380_ VGND VGND VPWR VPWR _06386_
+ sky130_fd_sc_hd__and2_1
XFILLER_28_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13785_ clknet_leaf_64_clk _00331_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10997_ sha256cu.m_pad_pars.m_size\[3\] sha256cu.m_pad_pars.block_512\[63\]\[3\]
+ _01919_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__mux2_1
X_12736_ sha256cu.m_pad_pars.block_512\[22\]\[5\] _06343_ VGND VGND VPWR VPWR _06349_
+ sky130_fd_sc_hd__and2_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12667_ _06312_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__clkbuf_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11618_ sha256cu.msg_scheduler.mreg_9\[1\] sha256cu.msg_scheduler.mreg_0\[1\] VGND
+ VGND VPWR VPWR _05450_ sky130_fd_sc_hd__or2_1
X_14406_ clknet_leaf_77_clk _00920_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[22\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12598_ sha256cu.m_pad_pars.block_512\[14\]\[4\] _06271_ VGND VGND VPWR VPWR _06276_
+ sky130_fd_sc_hd__and2_1
XFILLER_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14337_ clknet_leaf_105_clk _00851_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.counter_iteration\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11549_ sha256cu.data_in_padd\[30\] _01980_ _01987_ _05385_ VGND VGND VPWR VPWR _00893_
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14268_ clknet_leaf_19_clk _00814_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14199_ clknet_leaf_28_clk _00745_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_13219_ _06606_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__clkbuf_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _03237_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__nand2_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ _02113_ _02330_ _02331_ _02332_ sha256cu.m_out_digest.a_in\[8\] VGND VGND
+ VPWR VPWR _00103_ sky130_fd_sc_hd__a32o_1
X_08691_ sha256cu.iter_processing.w\[0\] _02020_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__nand2_1
X_07642_ _02262_ _02263_ _02264_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__and3_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07573_ sha256cu.m_out_digest.a_in\[18\] VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__clkbuf_4
X_09312_ _03789_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__nor2_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09243_ _03612_ _03720_ _03721_ _03724_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__o31a_2
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09174_ _03643_ _03627_ _03656_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__or3_1
X_08125_ _02705_ _02724_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__a21bo_1
XFILLER_147_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08056_ sha256cu.iter_processing.w\[17\] _02640_ _02667_ VGND VGND VPWR VPWR _02668_
+ sky130_fd_sc_hd__a21o_1
XFILLER_89_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07007_ _01644_ _01688_ _01689_ _01692_ _01629_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__o311a_1
XFILLER_1_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput116 hash[203] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput105 hash[194] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
Xinput127 hash[213] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08958_ sha256cu.m_out_digest.e_in\[10\] _02070_ _03449_ VGND VGND VPWR VPWR _00233_
+ sky130_fd_sc_hd__a21o_1
XFILLER_102_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput138 hash[223] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
Xinput149 hash[233] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
X_08889_ _03352_ _03353_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__or2_1
X_07909_ sha256cu.m_out_digest.e_in\[25\] _02524_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__xnor2_2
XFILLER_57_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10920_ _01956_ _04786_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__nand2_4
XFILLER_29_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10851_ sha256cu.m_pad_pars.add_out2\[5\] sha256cu.m_pad_pars.add_out2\[4\] VGND
+ VGND VPWR VPWR _04726_ sky130_fd_sc_hd__and2b_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10782_ sha256cu.msg_scheduler.mreg_12\[19\] _04679_ VGND VGND VPWR VPWR _04682_
+ sky130_fd_sc_hd__or2_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ clknet_leaf_85_clk _00116_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[21\]
+ sky130_fd_sc_hd__dfxtp_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ sha256cu.m_pad_pars.block_512\[10\]\[1\] _06232_ VGND VGND VPWR VPWR _06234_
+ sky130_fd_sc_hd__and2_1
XFILLER_40_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _06197_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11403_ _04819_ _05233_ _05246_ sha256cu.m_pad_pars.block_512\[37\]\[7\] VGND VGND
+ VPWR VPWR _05247_ sky130_fd_sc_hd__o22a_1
XFILLER_153_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12383_ sha256cu.m_pad_pars.block_512\[2\]\[0\] _06160_ VGND VGND VPWR VPWR _06161_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14122_ clknet_leaf_32_clk _00668_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11334_ sha256cu.m_pad_pars.block_512\[1\]\[2\] _05135_ _05151_ sha256cu.m_pad_pars.block_512\[49\]\[2\]
+ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__a22o_1
X_14053_ clknet_leaf_40_clk _00599_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11265_ _04702_ _04758_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__nor2_1
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10216_ sha256cu.msg_scheduler.mreg_3\[31\] _04354_ _04359_ _04357_ VGND VGND VPWR
+ VPWR _00587_ sky130_fd_sc_hd__o211a_1
X_13004_ sha256cu.m_pad_pars.block_512\[38\]\[2\] _06489_ VGND VGND VPWR VPWR _06492_
+ sky130_fd_sc_hd__and2_1
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11196_ sha256cu.m_pad_pars.block_512\[26\]\[4\] _04964_ _05014_ sha256cu.m_pad_pars.block_512\[18\]\[4\]
+ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a22o_1
X_10147_ sha256cu.msg_scheduler.mreg_3\[1\] _04315_ _04320_ _04318_ VGND VGND VPWR
+ VPWR _00557_ sky130_fd_sc_hd__o211a_1
XFILLER_121_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10078_ sha256cu.msg_scheduler.mreg_2\[4\] _04274_ _04280_ _04277_ VGND VGND VPWR
+ VPWR _00528_ sky130_fd_sc_hd__o211a_1
XFILLER_94_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14955_ clknet_leaf_105_clk _01469_ VGND VGND VPWR VPWR sha256cu.K\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13906_ clknet_leaf_96_clk _00452_ VGND VGND VPWR VPWR sha256cu.counter_iteration\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14886_ clknet_leaf_117_clk _01400_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13837_ clknet_leaf_18_clk _00383_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13768_ clknet_leaf_83_clk _00314_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_12719_ sha256cu.m_pad_pars.block_512\[21\]\[5\] _06334_ VGND VGND VPWR VPWR _06340_
+ sky130_fd_sc_hd__and2_1
X_13699_ clknet_leaf_85_clk _00245_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[22\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09930_ sha256cu.msg_scheduler.mreg_0\[4\] _04195_ _04196_ _04171_ VGND VGND VPWR
+ VPWR _00464_ sky130_fd_sc_hd__o211a_1
X_09861_ sha256cu.msg_scheduler.mreg_12\[16\] _04153_ _04154_ _04144_ VGND VGND VPWR
+ VPWR _00431_ sky130_fd_sc_hd__o211a_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _03307_ _03308_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__nor2_1
X_09792_ sha256cu.msg_scheduler.mreg_13\[19\] _04112_ _04114_ _04103_ VGND VGND VPWR
+ VPWR _00402_ sky130_fd_sc_hd__o211a_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ sha256cu.iter_processing.w\[3\] _02120_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__or2_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08674_ _02515_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__clkbuf_8
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07625_ sha256cu.K\[6\] _02248_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__xnor2_2
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07556_ _02104_ _02146_ _02145_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__o21a_1
X_07487_ _02113_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__buf_4
X_09226_ _03703_ _03707_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__nor2_1
XFILLER_10_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09157_ sha256cu.m_out_digest.e_in\[17\] _02040_ _03641_ _02068_ VGND VGND VPWR VPWR
+ _00240_ sky130_fd_sc_hd__a211o_1
X_09088_ _03540_ _03544_ _03538_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__o21a_1
X_08108_ _02676_ _02679_ _02718_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__o21a_1
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08039_ _02641_ _02651_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__xor2_1
XFILLER_116_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11050_ _04702_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__nor2_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10001_ _04116_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__buf_2
XFILLER_107_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14740_ clknet_leaf_5_clk _01254_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11952_ _05768_ _05769_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__or2b_1
XFILLER_44_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11883_ _05702_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__or2_2
XFILLER_45_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14671_ clknet_leaf_0_clk _01185_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[31\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10903_ _04748_ _01953_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__or2_2
X_13622_ clknet_leaf_63_clk _00168_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10834_ _04714_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
X_13553_ clknet_leaf_51_clk _00099_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_13_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10765_ _04580_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__buf_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12504_ sha256cu.m_pad_pars.block_512\[9\]\[1\] _06223_ VGND VGND VPWR VPWR _06225_
+ sky130_fd_sc_hd__and2_1
X_10696_ _04580_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__buf_2
XFILLER_9_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13484_ sha256cu.K\[20\] _06713_ _06718_ _00048_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__a22o_1
XFILLER_138_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12435_ _06188_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12366_ _01965_ _05244_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__nand2_2
XFILLER_153_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14105_ clknet_leaf_35_clk _00651_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11317_ sha256cu.m_pad_pars.block_512\[49\]\[0\] _05151_ _05158_ sha256cu.m_pad_pars.block_512\[21\]\[0\]
+ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a221o_1
X_12297_ sha256cu.msg_scheduler.mreg_1\[16\] sha256cu.msg_scheduler.mreg_1\[5\] VGND
+ VGND VPWR VPWR _06100_ sky130_fd_sc_hd__xor2_1
XFILLER_99_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14036_ clknet_leaf_39_clk _00582_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11248_ _04952_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__and2b_1
XFILLER_79_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11179_ _05032_ _05034_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__or3_1
XFILLER_68_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14938_ clknet_leaf_91_clk _01452_ VGND VGND VPWR VPWR sha256cu.K\[11\] sky130_fd_sc_hd__dfxtp_4
X_14869_ clknet_leaf_124_clk _01383_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07410_ _02039_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08390_ _02988_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__nor2_1
XFILLER_51_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07341_ _01982_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
X_07272_ sha256cu.m_pad_pars.block_512\[63\]\[0\] _01924_ VGND VGND VPWR VPWR _01925_
+ sky130_fd_sc_hd__and2_1
X_09011_ _03443_ _03447_ _03471_ _03500_ _03470_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a311oi_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09913_ _04185_ _04186_ _02007_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__and3b_1
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09844_ sha256cu.msg_scheduler.mreg_13\[9\] _04134_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__or2_1
XFILLER_59_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09775_ sha256cu.msg_scheduler.mreg_14\[12\] _04093_ VGND VGND VPWR VPWR _04105_
+ sky130_fd_sc_hd__or2_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06987_ _01602_ _01626_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__nor2_1
XFILLER_27_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ sha256cu.m_out_digest.h_in\[2\] sha256cu.m_out_digest.d_in\[2\] VGND VGND
+ VPWR VPWR _03226_ sky130_fd_sc_hd__nand2_1
XFILLER_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ sha256cu.m_out_digest.d_in\[3\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[3\]
+ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__o22a_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ sha256cu.m_out_digest.a_in\[28\] VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__buf_4
XFILLER_42_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08588_ sha256cu.m_out_digest.b_in\[10\] _02370_ _02110_ sha256cu.m_out_digest.a_in\[10\]
+ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__o22a_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07539_ sha256cu.m_out_digest.h_in\[4\] _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ sha256cu.msg_scheduler.mreg_8\[14\] _04540_ _04550_ _04543_ VGND VGND VPWR
+ VPWR _00730_ sky130_fd_sc_hd__o211a_1
X_10481_ sha256cu.msg_scheduler.mreg_7\[17\] _04500_ _04510_ _04503_ VGND VGND VPWR
+ VPWR _00701_ sky130_fd_sc_hd__o211a_1
XFILLER_136_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09209_ _03664_ _03666_ _03662_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__a21o_1
XFILLER_136_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12220_ _05983_ _06005_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nand2_1
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12151_ sha256cu.iter_processing.w\[23\] _05894_ _05960_ _05866_ VGND VGND VPWR VPWR
+ _00921_ sky130_fd_sc_hd__o211a_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12082_ _04043_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__clkbuf_4
X_11102_ _04701_ _04753_ _04960_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__o21a_1
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11033_ sha256cu.m_pad_pars.m_size\[6\] sha256cu.m_pad_pars.block_512\[63\]\[6\]
+ _01919_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__mux2_1
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12984_ _06481_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__clkbuf_1
X_11935_ _05750_ _05752_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__a21o_1
XFILLER_73_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14723_ clknet_leaf_99_clk _01237_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14654_ clknet_leaf_115_clk _01168_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11866_ sha256cu.iter_processing.w\[11\] _05666_ _05687_ _05640_ VGND VGND VPWR VPWR
+ _00909_ sky130_fd_sc_hd__o211a_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13605_ clknet_leaf_81_clk _00151_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11797_ sha256cu.msg_scheduler.mreg_9\[9\] sha256cu.msg_scheduler.mreg_0\[9\] VGND
+ VGND VPWR VPWR _05621_ sky130_fd_sc_hd__or2_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14585_ clknet_leaf_118_clk _01099_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10817_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__buf_4
X_10748_ sha256cu.msg_scheduler.mreg_12\[4\] _04653_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__or2_1
X_13536_ clknet_leaf_79_clk _00033_ VGND VGND VPWR VPWR state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13467_ sha256cu.K\[13\] _06726_ _06727_ _06743_ _06737_ VGND VGND VPWR VPWR _01454_
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10679_ sha256cu.msg_scheduler.mreg_11\[6\] _04614_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__or2_1
X_12418_ _06179_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13398_ _06700_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12349_ sha256cu.m_pad_pars.add_512_block\[6\] _06142_ _06143_ VGND VGND VPWR VPWR
+ _00936_ sky130_fd_sc_hd__o21ba_1
XFILLER_114_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14019_ clknet_leaf_56_clk _00565_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06910_ _01589_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07890_ _02443_ _02462_ _02506_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06841_ net10 net14 net13 net16 VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__or4_1
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09560_ sha256cu.m_out_digest.f_in\[3\] _03191_ _04026_ sha256cu.m_out_digest.e_in\[3\]
+ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__o22a_1
XFILLER_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09491_ _03961_ _03962_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__and2_1
X_08511_ _02272_ _02220_ _03109_ _03111_ _02258_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__a221o_1
X_08442_ sha256cu.m_out_digest.e_in\[7\] sha256cu.m_out_digest.e_in\[2\] VGND VGND
+ VPWR VPWR _03044_ sky130_fd_sc_hd__xnor2_4
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08373_ _02974_ _02976_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__xor2_1
X_07324_ _01962_ _01967_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__nor2_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07255_ net259 state\[3\] net257 VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__o21ba_1
X_07186_ _01650_ _01681_ _01851_ _01852_ _01629_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__o311a_1
XFILLER_145_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09827_ sha256cu.msg_scheduler.mreg_12\[1\] _04126_ _04135_ _04130_ VGND VGND VPWR
+ VPWR _00416_ sky130_fd_sc_hd__o211a_1
XFILLER_59_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09758_ sha256cu.msg_scheduler.mreg_13\[4\] _04086_ _04095_ _04090_ VGND VGND VPWR
+ VPWR _00387_ sky130_fd_sc_hd__o211a_1
XFILLER_27_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08709_ _03208_ _03209_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__xnor2_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ sha256cu.msg_scheduler.mreg_14\[6\] _04045_ _04056_ _04050_ VGND VGND VPWR
+ VPWR _00357_ sky130_fd_sc_hd__o211a_1
X_11720_ _05546_ _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nor2_1
XFILLER_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11651_ _05479_ _05480_ _05460_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__a21oi_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10602_ sha256cu.msg_scheduler.mreg_9\[5\] _04567_ _04579_ _04570_ VGND VGND VPWR
+ VPWR _00753_ sky130_fd_sc_hd__o211a_1
X_14370_ clknet_leaf_109_clk _00884_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11582_ _01935_ _05277_ _05413_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__a31o_1
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10533_ _04447_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__buf_2
X_13321_ _01923_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__buf_2
XFILLER_109_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10464_ sha256cu.msg_scheduler.mreg_8\[10\] _04494_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__or2_1
XFILLER_109_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13252_ sha256cu.m_pad_pars.block_512\[52\]\[6\] _06617_ VGND VGND VPWR VPWR _06624_
+ sky130_fd_sc_hd__and2_1
X_10395_ sha256cu.msg_scheduler.mreg_7\[12\] _04455_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__or2_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ sha256cu.msg_scheduler.mreg_9\[26\] sha256cu.msg_scheduler.mreg_0\[26\] VGND
+ VGND VPWR VPWR _06010_ sky130_fd_sc_hd__or2_1
X_13183_ sha256cu.m_pad_pars.block_512\[48\]\[6\] _06580_ VGND VGND VPWR VPWR _06587_
+ sky130_fd_sc_hd__and2_1
XFILLER_151_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12134_ sha256cu.msg_scheduler.mreg_1\[26\] sha256cu.msg_scheduler.mreg_1\[9\] VGND
+ VGND VPWR VPWR _05944_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12065_ sha256cu.msg_scheduler.mreg_14\[30\] _05877_ VGND VGND VPWR VPWR _05878_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_77_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11016_ sha256cu.m_pad_pars.block_512\[11\]\[4\] _04790_ _04831_ sha256cu.m_pad_pars.block_512\[19\]\[4\]
+ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__a22o_1
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12967_ _06472_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__clkbuf_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _05711_ _05715_ _05712_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__a21boi_1
XFILLER_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14706_ clknet_leaf_5_clk _01220_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12898_ _06435_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_360 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ sha256cu.msg_scheduler.mreg_1\[18\] sha256cu.msg_scheduler.mreg_1\[14\] VGND
+ VGND VPWR VPWR _05671_ sky130_fd_sc_hd__xnor2_1
XANTENNA_382 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14637_ clknet_leaf_12_clk _01151_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_393 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_371 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ clknet_leaf_14_clk _01082_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13519_ clknet_leaf_79_clk _00069_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dfxtp_2
X_14499_ clknet_leaf_103_clk _01013_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_07040_ _01602_ _01684_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__nand2_1
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08991_ _03479_ _03480_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07942_ _02520_ _02521_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__and2b_1
X_07873_ sha256cu.iter_processing.w\[13\] _02489_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09612_ _02515_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__clkbuf_4
X_06824_ _01518_ _01519_ _01520_ _01521_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__or4_1
X_09543_ _04011_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09474_ _03946_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__xor2_1
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08425_ _02988_ _02993_ _03027_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__o21ba_1
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08356_ _02128_ sha256cu.m_out_digest.a_in\[7\] VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07307_ sha256cu.m_pad_pars.add_512_block\[6\] _01950_ VGND VGND VPWR VPWR _01951_
+ sky130_fd_sc_hd__or2_1
XFILLER_149_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08287_ sha256cu.m_out_digest.h_in\[24\] _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07238_ _01849_ _01633_ _01611_ _01657_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__a211o_1
XFILLER_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07169_ _01790_ _01796_ _01837_ _01618_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__o22a_1
XFILLER_145_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10180_ sha256cu.msg_scheduler.mreg_4\[16\] _04335_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__or2_1
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13870_ clknet_leaf_20_clk _00416_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12821_ _06394_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ sha256cu.m_pad_pars.block_512\[23\]\[4\] _06353_ VGND VGND VPWR VPWR _06358_
+ sky130_fd_sc_hd__and2_1
X_11703_ sha256cu.msg_scheduler.mreg_9\[5\] sha256cu.msg_scheduler.mreg_0\[5\] VGND
+ VGND VPWR VPWR _05531_ sky130_fd_sc_hd__nand2_1
XFILLER_70_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ sha256cu.m_pad_pars.block_512\[19\]\[4\] _06316_ VGND VGND VPWR VPWR _06321_
+ sky130_fd_sc_hd__and2_1
XFILLER_43_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11634_ _05432_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__clkbuf_4
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ clknet_leaf_108_clk _00936_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_512_block\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_14353_ clknet_leaf_110_clk _00867_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11565_ _04815_ _04913_ _05302_ sha256cu.m_pad_pars.block_512\[36\]\[7\] VGND VGND
+ VPWR VPWR _05401_ sky130_fd_sc_hd__o22a_1
XFILLER_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10516_ sha256cu.msg_scheduler.mreg_9\[0\] _04520_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__or2_1
X_14284_ clknet_leaf_24_clk _00830_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11496_ sha256cu.m_pad_pars.block_512\[32\]\[2\] _05306_ _05318_ sha256cu.m_pad_pars.block_512\[8\]\[2\]
+ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__a221o_1
XFILLER_10_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13304_ _06651_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10447_ sha256cu.msg_scheduler.mreg_7\[2\] _04487_ _04491_ _04490_ VGND VGND VPWR
+ VPWR _00686_ sky130_fd_sc_hd__o211a_1
X_13235_ sha256cu.m_pad_pars.block_512\[51\]\[6\] _06608_ VGND VGND VPWR VPWR _06615_
+ sky130_fd_sc_hd__and2_1
X_10378_ sha256cu.msg_scheduler.mreg_6\[4\] _04448_ _04452_ _04451_ VGND VGND VPWR
+ VPWR _00656_ sky130_fd_sc_hd__o211a_1
X_13166_ sha256cu.m_pad_pars.block_512\[47\]\[6\] _06571_ VGND VGND VPWR VPWR _06578_
+ sky130_fd_sc_hd__and2_1
X_12117_ _05925_ _05926_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__or2_1
X_13097_ sha256cu.m_pad_pars.block_512\[43\]\[6\] _06534_ VGND VGND VPWR VPWR _06541_
+ sky130_fd_sc_hd__and2_1
X_12048_ _05838_ _05841_ _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13999_ clknet_leaf_56_clk _00545_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_190 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08210_ sha256cu.m_out_digest.b_in\[22\] _02026_ _02817_ VGND VGND VPWR VPWR _02818_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09190_ _03671_ _03672_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__nand2_1
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08141_ _02748_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__xnor2_2
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08072_ _02673_ _02683_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__xor2_1
XFILLER_146_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07023_ _01700_ _01705_ _01707_ _01652_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__o22a_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08974_ _03430_ _03435_ _03428_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__o21ba_1
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07925_ _02538_ _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07856_ _02409_ _02434_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__nor2_1
XFILLER_110_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07787_ _02401_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__xor2_1
X_06807_ net165 net169 net168 net171 VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__or4_1
XFILLER_44_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09526_ _03963_ _03970_ _03997_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__o21a_1
XFILLER_71_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09457_ _03929_ _03930_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__nand2_1
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08408_ _03005_ _03010_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__nand2_1
XFILLER_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09388_ _03863_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__and2b_1
X_08339_ _02925_ _02926_ _02942_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__and3_1
X_11350_ sha256cu.m_pad_pars.block_512\[49\]\[3\] _05151_ _05158_ sha256cu.m_pad_pars.block_512\[21\]\[3\]
+ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__a221o_1
XFILLER_153_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10301_ sha256cu.msg_scheduler.mreg_6\[4\] _04401_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__or2_1
XFILLER_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11281_ sha256cu.m_pad_pars.add_out1\[2\] _05125_ _05131_ sha256cu.m_pad_pars.add_out1\[3\]
+ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__and4b_2
X_13020_ _06500_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__clkbuf_1
X_10232_ sha256cu.msg_scheduler.mreg_4\[6\] _04367_ _04368_ _04357_ VGND VGND VPWR
+ VPWR _00594_ sky130_fd_sc_hd__o211a_1
XFILLER_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10163_ sha256cu.msg_scheduler.mreg_3\[8\] _04328_ _04329_ _04318_ VGND VGND VPWR
+ VPWR _00564_ sky130_fd_sc_hd__o211a_1
XFILLER_120_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10094_ sha256cu.msg_scheduler.mreg_3\[11\] _04282_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__or2_1
XFILLER_87_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13922_ clknet_leaf_44_clk _00468_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13853_ clknet_leaf_22_clk _00399_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12804_ _06385_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13784_ clknet_leaf_63_clk _00330_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10996_ sha256cu.data_in_padd\[2\] _04840_ _04852_ _04860_ _01974_ VGND VGND VPWR
+ VPWR _00865_ sky130_fd_sc_hd__o221a_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _06348_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__clkbuf_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12666_ sha256cu.m_pad_pars.block_512\[18\]\[4\] _06307_ VGND VGND VPWR VPWR _06312_
+ sky130_fd_sc_hd__and2_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ sha256cu.msg_scheduler.mreg_9\[1\] sha256cu.msg_scheduler.mreg_0\[1\] VGND
+ VGND VPWR VPWR _05449_ sky130_fd_sc_hd__nand2_1
X_12597_ _06275_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__clkbuf_1
X_14405_ clknet_leaf_76_clk _00919_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[21\]
+ sky130_fd_sc_hd__dfxtp_2
X_14336_ clknet_leaf_10_clk _00850_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.m_size\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11548_ _05377_ _05379_ _05384_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__or3_2
X_14267_ clknet_leaf_19_clk _00813_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11479_ sha256cu.m_pad_pars.block_512\[4\]\[0\] _05313_ _05314_ sha256cu.m_pad_pars.block_512\[0\]\[0\]
+ _05321_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__a221o_1
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14198_ clknet_leaf_28_clk _00744_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13218_ sha256cu.m_pad_pars.block_512\[50\]\[6\] _06599_ VGND VGND VPWR VPWR _06606_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13149_ sha256cu.m_pad_pars.block_512\[46\]\[6\] _06562_ VGND VGND VPWR VPWR _06569_
+ sky130_fd_sc_hd__and2_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07710_ _02065_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__buf_4
XFILLER_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08690_ sha256cu.m_out_digest.d_in\[31\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[31\]
+ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__o22a_1
XFILLER_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07641_ sha256cu.m_out_digest.g_in\[7\] sha256cu.m_out_digest.f_in\[7\] sha256cu.m_out_digest.e_in\[7\]
+ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__mux2_1
XFILLER_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07572_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__inv_2
XFILLER_81_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09311_ _02811_ _03757_ _03758_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a21boi_1
XFILLER_22_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09242_ _03690_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__nor2_1
X_09173_ _03643_ _03627_ _03656_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__o21ai_1
X_08124_ _02723_ _02721_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__or2b_1
XFILLER_147_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08055_ _02638_ _02639_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__and2b_1
XFILLER_143_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07006_ _01690_ _01603_ _01612_ _01691_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__a31o_1
XFILLER_1_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput106 hash[195] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
XFILLER_102_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput117 hash[204] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
X_08957_ _03443_ _03445_ _03447_ _03448_ _02113_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__o311a_1
XFILLER_130_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput139 hash[224] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput128 hash[214] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08888_ _03376_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__xor2_1
X_07908_ sha256cu.m_out_digest.e_in\[20\] sha256cu.m_out_digest.e_in\[7\] VGND VGND
+ VPWR VPWR _02524_ sky130_fd_sc_hd__xnor2_1
X_07839_ _02418_ _02421_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__o21a_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10850_ sha256cu.m_pad_pars.add_out2\[5\] VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10781_ sha256cu.msg_scheduler.mreg_11\[18\] _04672_ _04681_ _04675_ VGND VGND VPWR
+ VPWR _00830_ sky130_fd_sc_hd__o211a_1
X_09509_ _03951_ _03954_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__a21oi_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _06233_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ sha256cu.m_pad_pars.block_512\[6\]\[0\] _06196_ VGND VGND VPWR VPWR _06197_
+ sky130_fd_sc_hd__and2_1
XFILLER_40_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11402_ _04792_ _04969_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__nor2_1
X_14121_ clknet_leaf_32_clk _00667_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12382_ _01965_ _04998_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__nand2_2
XANTENNA_90 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11333_ sha256cu.m_pad_pars.block_512\[13\]\[2\] _05128_ _05132_ sha256cu.m_pad_pars.block_512\[41\]\[2\]
+ _05181_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__a221o_1
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14052_ clknet_leaf_40_clk _00598_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11264_ _04727_ _05102_ _05106_ _05115_ _01969_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__a2111o_1
X_10215_ sha256cu.msg_scheduler.mreg_4\[31\] _04348_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__or2_1
XFILLER_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13003_ _06491_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11195_ sha256cu.data_in_padd\[11\] _04840_ _05047_ _05050_ _05040_ VGND VGND VPWR
+ VPWR _00874_ sky130_fd_sc_hd__o221a_1
XFILLER_0_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10146_ sha256cu.msg_scheduler.mreg_4\[1\] _04308_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__or2_1
XFILLER_121_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10077_ sha256cu.msg_scheduler.mreg_3\[4\] _04268_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__or2_1
X_14954_ clknet_leaf_89_clk _01468_ VGND VGND VPWR VPWR sha256cu.K\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13905_ clknet_leaf_105_clk _00451_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.counter_iteration\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_36_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14885_ clknet_leaf_99_clk _01399_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13836_ clknet_leaf_76_clk _00382_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[31\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13767_ clknet_leaf_82_clk _00313_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10979_ sha256cu.m_pad_pars.block_512\[27\]\[1\] _04757_ _04828_ sha256cu.m_pad_pars.block_512\[23\]\[1\]
+ _04844_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__a221o_1
XFILLER_16_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12718_ _06339_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_1
X_13698_ clknet_leaf_84_clk _00244_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[21\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12649_ sha256cu.m_pad_pars.block_512\[17\]\[4\] _06298_ VGND VGND VPWR VPWR _06303_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14319_ clknet_leaf_91_clk _00013_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09860_ sha256cu.msg_scheduler.mreg_13\[16\] _04147_ VGND VGND VPWR VPWR _04154_
+ sky130_fd_sc_hd__or2_1
XFILLER_98_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _03290_ _03280_ _03306_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__and3_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09791_ sha256cu.msg_scheduler.mreg_14\[19\] _04106_ VGND VGND VPWR VPWR _04114_
+ sky130_fd_sc_hd__or2_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08742_ sha256cu.iter_processing.w\[3\] _02120_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__nand2_1
XFILLER_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08673_ sha256cu.m_out_digest.d_in\[16\] _03187_ _03190_ sha256cu.m_out_digest.c_in\[16\]
+ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__o22a_1
XFILLER_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07624_ _02245_ _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__xor2_2
XFILLER_93_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ _02178_ _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__xor2_1
X_07486_ _02112_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__buf_4
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09225_ sha256cu.K\[20\] _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09156_ _02069_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__nor2_1
XFILLER_147_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09087_ _03568_ _03573_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__xor2_1
X_08107_ sha256cu.m_out_digest.h_in\[18\] _02678_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_110_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_16
X_08038_ _02648_ _02650_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10000_ sha256cu.msg_scheduler.mreg_2\[3\] _04228_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__or2_1
XFILLER_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09989_ sha256cu.msg_scheduler.mreg_1\[30\] _04228_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__or2_1
XFILLER_103_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11951_ _05738_ _05743_ _05767_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__a21o_1
XFILLER_57_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11882_ _05677_ _05679_ _05675_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__a21oi_1
X_14670_ clknet_leaf_110_clk _01184_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10902_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__buf_4
XFILLER_45_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13621_ clknet_leaf_61_clk _00167_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10833_ sha256cu.m_pad_pars.m_size\[9\] _01994_ _04700_ VGND VGND VPWR VPWR _04714_
+ sky130_fd_sc_hd__and3_1
X_13552_ clknet_leaf_51_clk _00098_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[3\]
+ sky130_fd_sc_hd__dfxtp_4
X_10764_ sha256cu.msg_scheduler.mreg_11\[11\] _04659_ _04671_ _04662_ VGND VGND VPWR
+ VPWR _00823_ sky130_fd_sc_hd__o211a_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12503_ _06224_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
X_10695_ sha256cu.msg_scheduler.mreg_10\[13\] _04620_ _04632_ _04623_ VGND VGND VPWR
+ VPWR _00793_ sky130_fd_sc_hd__o211a_1
XFILLER_9_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13483_ sha256cu.K\[19\] _06726_ _06727_ _06753_ _06737_ VGND VGND VPWR VPWR _01460_
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12434_ sha256cu.m_pad_pars.block_512\[5\]\[0\] _06187_ VGND VGND VPWR VPWR _06188_
+ sky130_fd_sc_hd__and2_1
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_101_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_16
X_12365_ _01984_ _01942_ _04775_ sha256cu.m_pad_pars.block_512\[0\]\[7\] VGND VGND
+ VPWR VPWR _00944_ sky130_fd_sc_hd__a31o_1
XFILLER_153_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14104_ clknet_leaf_36_clk _00650_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11316_ sha256cu.m_pad_pars.block_512\[5\]\[0\] _05160_ _05161_ sha256cu.m_pad_pars.block_512\[53\]\[0\]
+ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a221o_1
X_14035_ clknet_leaf_39_clk _00581_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12296_ _06097_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__nand2_1
XFILLER_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11247_ sha256cu.m_pad_pars.block_512\[6\]\[7\] _04955_ _04954_ _04933_ VGND VGND
+ VPWR VPWR _05099_ sky130_fd_sc_hd__o22a_1
XFILLER_122_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11178_ sha256cu.m_pad_pars.block_512\[30\]\[2\] _05009_ _04977_ sha256cu.m_pad_pars.block_512\[46\]\[2\]
+ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__a22o_1
X_10129_ sha256cu.msg_scheduler.mreg_3\[26\] _04308_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__or2_1
XFILLER_121_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14937_ clknet_leaf_91_clk _01451_ VGND VGND VPWR VPWR sha256cu.K\[10\] sky130_fd_sc_hd__dfxtp_4
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14868_ clknet_leaf_1_clk _01382_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13819_ clknet_leaf_47_clk _00365_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_07340_ _01975_ _01978_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__and3_1
X_14799_ clknet_leaf_0_clk _01313_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09010_ _03441_ _03469_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__nor2_1
X_07271_ _01923_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__clkbuf_2
XFILLER_31_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09912_ sha256cu.msg_scheduler.counter_iteration\[4\] _04181_ sha256cu.msg_scheduler.counter_iteration\[5\]
+ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a21o_1
XFILLER_98_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09843_ sha256cu.msg_scheduler.mreg_12\[8\] _04140_ _04143_ _04144_ VGND VGND VPWR
+ VPWR _00423_ sky130_fd_sc_hd__o211a_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09774_ sha256cu.msg_scheduler.mreg_13\[11\] _04099_ _04104_ _04103_ VGND VGND VPWR
+ VPWR _00394_ sky130_fd_sc_hd__o211a_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _01578_ _01606_ _01589_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__and3_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _02071_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _02515_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__buf_4
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ sha256cu.m_out_digest.b_in\[9\] _02370_ _02110_ sha256cu.m_out_digest.a_in\[9\]
+ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__o22a_1
X_07607_ _02230_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__inv_2
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07538_ _02161_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07469_ _02032_ _02060_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__or2_1
X_10480_ sha256cu.msg_scheduler.mreg_8\[17\] _04507_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__or2_1
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09208_ _03689_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__nor2_1
XFILLER_10_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09139_ sha256cu.iter_processing.w\[17\] _02639_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__and2_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12150_ _05442_ _05958_ _05959_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__a21o_1
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11101_ _04749_ _04953_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__or2_4
XFILLER_150_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12081_ sha256cu.iter_processing.w\[20\] _05666_ _05893_ _05866_ VGND VGND VPWR VPWR
+ _00918_ sky130_fd_sc_hd__o211a_1
XFILLER_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11032_ _01971_ _04892_ _04893_ _04709_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__o211a_1
XFILLER_89_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12983_ sha256cu.m_pad_pars.block_512\[37\]\[0\] _06480_ VGND VGND VPWR VPWR _06481_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11934_ sha256cu.data_in_padd\[14\] _05447_ _04692_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__a21o_1
XFILLER_73_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14722_ clknet_leaf_101_clk _01236_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14653_ clknet_leaf_123_clk _01167_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11865_ sha256cu.data_in_padd\[11\] _05667_ _05686_ _05463_ VGND VGND VPWR VPWR _05687_
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13604_ clknet_leaf_86_clk _00150_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11796_ _05612_ _05613_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__or2_1
XFILLER_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10816_ sha256cu.byte_rdy _01945_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__or2_4
X_14584_ clknet_leaf_120_clk _01098_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10747_ sha256cu.msg_scheduler.mreg_11\[3\] _04659_ _04661_ _04662_ VGND VGND VPWR
+ VPWR _00815_ sky130_fd_sc_hd__o211a_1
X_13535_ clknet_leaf_109_clk _00032_ VGND VGND VPWR VPWR state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10678_ sha256cu.msg_scheduler.mreg_10\[5\] _04620_ _04622_ _04623_ VGND VGND VPWR
+ VPWR _00785_ sky130_fd_sc_hd__o211a_1
X_13466_ _04188_ _00040_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__and2b_1
X_12417_ sha256cu.m_pad_pars.block_512\[4\]\[0\] _06178_ VGND VGND VPWR VPWR _06179_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13397_ sha256cu.m_pad_pars.block_512\[61\]\[3\] _06693_ VGND VGND VPWR VPWR _06700_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ sha256cu.m_pad_pars.add_512_block\[6\] _06142_ _02002_ VGND VGND VPWR VPWR
+ _06143_ sky130_fd_sc_hd__a21o_1
X_12279_ _06081_ _06082_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__xor2_1
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14018_ clknet_leaf_56_clk _00564_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06840_ _01522_ _01527_ _01532_ _01537_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__or4_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09490_ _03961_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__nor2_1
X_08510_ _02069_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__nor2_1
XFILLER_36_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08441_ sha256cu.m_out_digest.h_in\[28\] _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08372_ _02936_ _02941_ _02975_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__a21bo_1
XFILLER_149_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07323_ sha256cu.m_pad_pars.add_out1\[2\] _01963_ _01966_ VGND VGND VPWR VPWR _01967_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_32_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07254_ _01909_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07185_ _01637_ _01603_ _01701_ _01775_ _01620_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__a311o_1
XFILLER_117_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09826_ sha256cu.msg_scheduler.mreg_13\[1\] _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__or2_1
X_09757_ sha256cu.msg_scheduler.mreg_14\[4\] _04093_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__or2_1
XFILLER_74_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06969_ _01607_ _01605_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__nor2_2
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _02024_ _03199_ _03198_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__a21boi_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ sha256cu.iter_processing.w\[6\] _04054_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__or2_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08639_ sha256cu.m_out_digest.c_in\[19\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[19\]
+ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o22a_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11650_ _05460_ _05479_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__and3_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ sha256cu.msg_scheduler.mreg_10\[5\] _04574_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__or2_1
X_11581_ sha256cu.m_pad_pars.add_out0\[5\] sha256cu.m_pad_pars.add_out0\[4\] _05293_
+ _05415_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__a41o_1
X_10532_ sha256cu.msg_scheduler.mreg_8\[7\] _04526_ _04539_ _04530_ VGND VGND VPWR
+ VPWR _00723_ sky130_fd_sc_hd__o211a_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13320_ _06659_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10463_ _04447_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13251_ _06623_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
X_10394_ _04447_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__buf_2
XFILLER_136_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12202_ sha256cu.iter_processing.w\[25\] _05894_ _06009_ _05866_ VGND VGND VPWR VPWR
+ _00923_ sky130_fd_sc_hd__o211a_1
X_13182_ _06586_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__clkbuf_1
X_12133_ _05941_ _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__nand2_1
XFILLER_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12064_ sha256cu.msg_scheduler.mreg_14\[7\] sha256cu.msg_scheduler.mreg_14\[5\] VGND
+ VGND VPWR VPWR _05877_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11015_ sha256cu.m_pad_pars.block_512\[23\]\[4\] _04828_ _04818_ sha256cu.m_pad_pars.block_512\[35\]\[4\]
+ _04877_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__a221o_1
XFILLER_64_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12966_ sha256cu.m_pad_pars.block_512\[36\]\[0\] _06471_ VGND VGND VPWR VPWR _06472_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14705_ clknet_leaf_1_clk _01219_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_350 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _05733_ _05735_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__xor2_1
X_12897_ sha256cu.m_pad_pars.block_512\[32\]\[0\] _06434_ VGND VGND VPWR VPWR _06435_
+ sky130_fd_sc_hd__and2_1
XANTENNA_361 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_394 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _05668_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__nand2_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_372 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14636_ clknet_leaf_21_clk _01150_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_383 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567_ clknet_leaf_16_clk _01081_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11779_ _05570_ _05574_ _05571_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__a21boi_1
X_13518_ clknet_leaf_108_clk _00068_ VGND VGND VPWR VPWR sha256cu.byte_stop sky130_fd_sc_hd__dfxtp_1
XFILLER_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14498_ clknet_leaf_105_clk _01012_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13449_ sha256cu.K\[6\] _06714_ _06719_ _00064_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__a22o_1
XFILLER_142_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08990_ _02417_ _03454_ _03453_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__a21oi_1
X_07941_ sha256cu.K\[14\] _02541_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__nand2_1
X_07872_ _02487_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__xnor2_1
X_09611_ sha256cu.m_out_digest.g_in\[14\] _04032_ _04034_ sha256cu.m_out_digest.f_in\[14\]
+ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__o22a_1
XFILLER_95_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06823_ net90 net93 net92 net95 VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__or4_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09542_ _03159_ _04012_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09473_ sha256cu.K\[27\] _03907_ _03909_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_90_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_52_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08424_ _02986_ _02987_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__nor2_1
XFILLER_52_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08355_ _02945_ _02947_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__nor2_1
XFILLER_149_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07306_ sha256cu.m_pad_pars.add_512_block\[5\] sha256cu.m_pad_pars.add_512_block\[4\]
+ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__nand2_2
X_08286_ _02161_ _02891_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07237_ _01889_ _01891_ _01896_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07168_ _01657_ _01646_ _01611_ _01661_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__o31a_1
XFILLER_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07099_ _01654_ _01653_ _01776_ _01652_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__a211o_1
XFILLER_115_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09809_ sha256cu.msg_scheduler.mreg_13\[26\] _04112_ _04124_ _04117_ VGND VGND VPWR
+ VPWR _00409_ sky130_fd_sc_hd__o211a_1
XFILLER_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12820_ sha256cu.m_pad_pars.block_512\[27\]\[4\] _06389_ VGND VGND VPWR VPWR _06394_
+ sky130_fd_sc_hd__and2_1
XFILLER_28_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12751_ _06357_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11702_ sha256cu.msg_scheduler.mreg_9\[5\] sha256cu.msg_scheduler.mreg_0\[5\] VGND
+ VGND VPWR VPWR _05530_ sky130_fd_sc_hd__or2_1
XFILLER_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12682_ _06320_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11633_ sha256cu.iter_processing.w\[1\] _05430_ _05464_ _05335_ VGND VGND VPWR VPWR
+ _00899_ sky130_fd_sc_hd__o211a_1
XFILLER_70_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ clknet_leaf_112_clk _00935_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_512_block\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14352_ clknet_leaf_14_clk _00866_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11564_ _04801_ _05316_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__a21oi_1
X_10515_ sha256cu.msg_scheduler.mreg_7\[31\] _04526_ _04528_ _04530_ VGND VGND VPWR
+ VPWR _00715_ sky130_fd_sc_hd__o211a_1
XFILLER_109_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14283_ clknet_leaf_25_clk _00829_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11495_ sha256cu.m_pad_pars.block_512\[24\]\[2\] _05279_ _05298_ sha256cu.m_pad_pars.block_512\[44\]\[2\]
+ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__a22o_1
XFILLER_10_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13303_ sha256cu.m_pad_pars.block_512\[55\]\[6\] _06644_ VGND VGND VPWR VPWR _06651_
+ sky130_fd_sc_hd__and2_1
X_10446_ sha256cu.msg_scheduler.mreg_8\[2\] _04481_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__or2_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13234_ _06614_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10377_ sha256cu.msg_scheduler.mreg_7\[4\] _04441_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__or2_1
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13165_ _06577_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12116_ _05925_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__nand2_1
X_13096_ _06540_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__clkbuf_1
X_12047_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__inv_2
XFILLER_77_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13998_ clknet_leaf_56_clk _00544_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12949_ sha256cu.m_pad_pars.block_512\[35\]\[0\] _06462_ VGND VGND VPWR VPWR _06463_
+ sky130_fd_sc_hd__and2_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_72_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_180 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14619_ clknet_leaf_126_clk _01133_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08140_ _02713_ _02716_ _02749_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__o21a_1
X_08071_ _02680_ _02682_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__xnor2_1
X_07022_ _01690_ _01640_ _01706_ _01595_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__a31o_1
XFILLER_103_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08973_ _03462_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nor2_1
XFILLER_115_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07924_ _02485_ _02504_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__a21bo_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07855_ _02409_ _02434_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__nand2_1
XFILLER_84_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07786_ _02329_ _02403_ _02405_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__o21ba_1
X_06806_ Hash_Digest net1 VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__xor2_1
XFILLER_71_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09525_ _03992_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__xor2_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
X_09456_ sha256cu.m_out_digest.h_in\[28\] sha256cu.m_out_digest.d_in\[28\] VGND VGND
+ VPWR VPWR _03930_ sky130_fd_sc_hd__or2_1
XFILLER_40_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08407_ sha256cu.iter_processing.w\[27\] _03009_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__xor2_1
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09387_ _03826_ _03842_ _03862_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__a21o_1
XFILLER_40_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08338_ _02925_ _02926_ _02942_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08269_ _02874_ _02875_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10300_ _04314_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__buf_2
X_11280_ _04913_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__or2_1
X_10231_ sha256cu.msg_scheduler.mreg_5\[6\] _04361_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__or2_1
XFILLER_106_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10162_ sha256cu.msg_scheduler.mreg_4\[8\] _04322_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__or2_1
XFILLER_126_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10093_ sha256cu.msg_scheduler.mreg_2\[10\] _04288_ _04289_ _04277_ VGND VGND VPWR
+ VPWR _00534_ sky130_fd_sc_hd__o211a_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13921_ clknet_leaf_44_clk _00467_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13852_ clknet_leaf_21_clk _00398_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13783_ clknet_leaf_63_clk _00329_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12803_ sha256cu.m_pad_pars.block_512\[26\]\[4\] _06380_ VGND VGND VPWR VPWR _06385_
+ sky130_fd_sc_hd__and2_1
XFILLER_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_90_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12734_ sha256cu.m_pad_pars.block_512\[22\]\[4\] _06343_ VGND VGND VPWR VPWR _06348_
+ sky130_fd_sc_hd__and2_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10995_ sha256cu.m_pad_pars.block_512\[51\]\[2\] _04826_ _04853_ _04859_ VGND VGND
+ VPWR VPWR _04860_ sky130_fd_sc_hd__a211o_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _06311_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__clkbuf_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__buf_2
X_14404_ clknet_leaf_76_clk _00918_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[20\]
+ sky130_fd_sc_hd__dfxtp_4
X_12596_ sha256cu.m_pad_pars.block_512\[14\]\[3\] _06271_ VGND VGND VPWR VPWR _06275_
+ sky130_fd_sc_hd__and2_1
X_14335_ clknet_leaf_10_clk _00849_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.m_size\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11547_ sha256cu.m_pad_pars.block_512\[52\]\[6\] _05310_ _05380_ _05383_ VGND VGND
+ VPWR VPWR _05384_ sky130_fd_sc_hd__a211o_1
XFILLER_11_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14266_ clknet_leaf_19_clk _00812_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11478_ sha256cu.m_pad_pars.block_512\[8\]\[0\] _05318_ _05320_ sha256cu.m_pad_pars.block_512\[40\]\[0\]
+ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__a22o_1
X_14197_ clknet_leaf_29_clk _00743_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10429_ _04414_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__clkbuf_2
X_13217_ _06605_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13148_ _06568_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__clkbuf_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13079_ _06531_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__clkbuf_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07640_ sha256cu.m_out_digest.b_in\[7\] sha256cu.m_out_digest.a_in\[7\] sha256cu.m_out_digest.c_in\[7\]
+ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__a21o_1
XFILLER_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07571_ sha256cu.m_out_digest.e_in\[30\] _02195_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__xnor2_4
XFILLER_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_81_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09310_ _02851_ _03788_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__xor2_1
XFILLER_46_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09241_ _03664_ _03665_ _03691_ _03722_ _03662_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__a32o_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09172_ _03654_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__nor2_1
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08123_ _02332_ _02731_ _02733_ _01984_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__o211ai_1
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ _02636_ _02655_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__a21bo_1
XFILLER_135_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07005_ _01583_ _01597_ _01689_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__or3_1
XFILLER_134_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput118 hash[205] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_4
Xinput107 hash[196] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
X_08956_ _03445_ _03447_ _03443_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__o21ai_1
Xinput129 hash[215] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_08887_ _03377_ _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__xnor2_1
X_07907_ sha256cu.iter_processing.w\[14\] _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__xnor2_1
X_07838_ sha256cu.m_out_digest.h_in\[11\] _02420_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__nand2_1
XFILLER_84_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07769_ _02386_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_36_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
X_09508_ _03979_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__nor2_1
X_10780_ sha256cu.msg_scheduler.mreg_12\[18\] _04679_ VGND VGND VPWR VPWR _04681_
+ sky130_fd_sc_hd__or2_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _03912_ _03913_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__nor2_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _01965_ _04956_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__nand2_2
XFILLER_12_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11401_ sha256cu.m_pad_pars.block_512\[1\]\[7\] _05244_ _05134_ _05127_ VGND VGND
+ VPWR VPWR _05245_ sky130_fd_sc_hd__o211a_1
XFILLER_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14120_ clknet_leaf_32_clk _00666_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_80 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _02000_ _05244_ sha256cu.m_pad_pars.block_512\[1\]\[7\] VGND VGND VPWR VPWR
+ _00952_ sky130_fd_sc_hd__a21o_1
XFILLER_153_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11332_ sha256cu.m_pad_pars.block_512\[45\]\[2\] _05126_ VGND VGND VPWR VPWR _05181_
+ sky130_fd_sc_hd__and2_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14051_ clknet_leaf_40_clk _00597_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11263_ _04726_ _04990_ _05108_ _05110_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__a311o_1
XFILLER_4_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10214_ sha256cu.msg_scheduler.mreg_3\[30\] _04354_ _04358_ _04357_ VGND VGND VPWR
+ VPWR _00586_ sky130_fd_sc_hd__o211a_1
XFILLER_121_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11194_ sha256cu.m_pad_pars.block_512\[22\]\[3\] _05013_ _05049_ _01970_ VGND VGND
+ VPWR VPWR _05050_ sky130_fd_sc_hd__a211o_1
X_13002_ sha256cu.m_pad_pars.block_512\[38\]\[1\] _06489_ VGND VGND VPWR VPWR _06491_
+ sky130_fd_sc_hd__and2_1
XFILLER_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10145_ sha256cu.msg_scheduler.mreg_3\[0\] _04315_ _04319_ _04318_ VGND VGND VPWR
+ VPWR _00556_ sky130_fd_sc_hd__o211a_1
XFILLER_153_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10076_ sha256cu.msg_scheduler.mreg_2\[3\] _04274_ _04279_ _04277_ VGND VGND VPWR
+ VPWR _00527_ sky130_fd_sc_hd__o211a_1
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14953_ clknet_leaf_90_clk _01467_ VGND VGND VPWR VPWR sha256cu.K\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14884_ clknet_leaf_100_clk _01398_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13904_ clknet_leaf_105_clk _00450_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.counter_iteration\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_75_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13835_ clknet_leaf_76_clk _00381_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[30\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_63_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13766_ clknet_leaf_81_clk _00312_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10978_ sha256cu.m_pad_pars.block_512\[11\]\[1\] _04790_ _04831_ sha256cu.m_pad_pars.block_512\[19\]\[1\]
+ _04843_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a221o_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13697_ clknet_leaf_83_clk _00243_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[20\]
+ sky130_fd_sc_hd__dfxtp_4
X_12717_ sha256cu.m_pad_pars.block_512\[21\]\[4\] _06334_ VGND VGND VPWR VPWR _06339_
+ sky130_fd_sc_hd__and2_1
X_12648_ _06302_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12579_ _06265_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14318_ clknet_leaf_93_clk _00012_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14249_ clknet_leaf_26_clk _00795_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _03290_ _03280_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__a21oi_2
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09790_ sha256cu.msg_scheduler.mreg_13\[18\] _04112_ _04113_ _04103_ VGND VGND VPWR
+ VPWR _00401_ sky130_fd_sc_hd__o211a_1
XFILLER_58_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _02071_ _03224_ _03222_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__o21ai_2
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08672_ _02109_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__buf_4
XFILLER_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07623_ _02187_ _02209_ _02246_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__a21boi_2
XFILLER_54_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07554_ sha256cu.K\[3\] _02143_ _02179_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__a21oi_2
X_07485_ _02111_ _02037_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__nor2_4
X_09224_ _03704_ _03705_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__nor2_1
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09155_ _03637_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09086_ sha256cu.K\[15\] _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__xor2_1
X_08106_ _02713_ _02716_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08037_ _02600_ _02603_ _02649_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__o21a_1
XFILLER_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09988_ sha256cu.msg_scheduler.mreg_0\[29\] _04221_ _04229_ _04224_ VGND VGND VPWR
+ VPWR _00489_ sky130_fd_sc_hd__o211a_1
XFILLER_88_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08939_ sha256cu.K\[10\] VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__inv_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11950_ _05738_ _05743_ _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__and3_1
X_10901_ _01944_ _04699_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__nand2_4
XFILLER_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11881_ _05700_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__nand2_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13620_ clknet_leaf_59_clk _00166_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10832_ sha256cu.m_pad_pars.add_512_block\[5\] _04700_ _04713_ _04709_ VGND VGND
+ VPWR VPWR _00849_ sky130_fd_sc_hd__o211a_1
XFILLER_25_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13551_ clknet_leaf_73_clk _00097_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[2\]
+ sky130_fd_sc_hd__dfxtp_4
X_10763_ sha256cu.msg_scheduler.mreg_12\[11\] _04666_ VGND VGND VPWR VPWR _04671_
+ sky130_fd_sc_hd__or2_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12502_ sha256cu.m_pad_pars.block_512\[9\]\[0\] _06223_ VGND VGND VPWR VPWR _06224_
+ sky130_fd_sc_hd__and2_1
XFILLER_139_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10694_ sha256cu.msg_scheduler.mreg_11\[13\] _04627_ VGND VGND VPWR VPWR _04632_
+ sky130_fd_sc_hd__or2_1
X_13482_ sha256cu.counter_iteration\[6\] _00046_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__and2b_1
X_12433_ _01986_ _04933_ _05159_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__or3_2
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12364_ _06151_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14103_ clknet_leaf_35_clk _00649_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11315_ _05024_ _05164_ _05165_ sha256cu.m_pad_pars.block_512\[37\]\[0\] VGND VGND
+ VPWR VPWR _05166_ sky130_fd_sc_hd__a22o_1
XFILLER_153_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14034_ clknet_leaf_40_clk _00580_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_12295_ sha256cu.msg_scheduler.mreg_9\[30\] sha256cu.msg_scheduler.mreg_0\[30\] VGND
+ VGND VPWR VPWR _06098_ sky130_fd_sc_hd__nand2_1
XFILLER_99_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11246_ _04987_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__and2b_1
XFILLER_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11177_ sha256cu.m_pad_pars.block_512\[10\]\[2\] _04963_ _05001_ sha256cu.m_pad_pars.block_512\[42\]\[2\]
+ _05033_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__a221o_1
X_10128_ sha256cu.msg_scheduler.mreg_2\[25\] _04301_ _04309_ _04304_ VGND VGND VPWR
+ VPWR _00549_ sky130_fd_sc_hd__o211a_1
X_10059_ sha256cu.msg_scheduler.mreg_2\[28\] _04268_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__or2_1
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14936_ clknet_leaf_91_clk _01450_ VGND VGND VPWR VPWR sha256cu.K\[9\] sky130_fd_sc_hd__dfxtp_4
XFILLER_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14867_ clknet_leaf_1_clk _01381_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13818_ clknet_leaf_48_clk _00364_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_14798_ clknet_leaf_111_clk _01312_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13749_ clknet_leaf_65_clk _00295_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07270_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
X_09911_ sha256cu.msg_scheduler.counter_iteration\[5\] sha256cu.msg_scheduler.counter_iteration\[4\]
+ _04181_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__and3_1
XFILLER_132_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09842_ _04116_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__buf_2
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09773_ sha256cu.msg_scheduler.mreg_14\[11\] _04093_ VGND VGND VPWR VPWR _04104_
+ sky130_fd_sc_hd__or2_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _03222_ _03223_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__nand2_1
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _01608_ _01623_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__or2_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ sha256cu.m_out_digest.d_in\[2\] _03184_ _03182_ sha256cu.m_out_digest.c_in\[2\]
+ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__a22o_1
XFILLER_66_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08586_ sha256cu.m_out_digest.b_in\[8\] _03031_ _02114_ sha256cu.m_out_digest.a_in\[8\]
+ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__a22o_1
X_07606_ sha256cu.m_out_digest.e_in\[31\] _02229_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__xnor2_2
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07537_ _02162_ sha256cu.m_out_digest.a_in\[6\] VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07468_ _02072_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09207_ _03657_ _03669_ _03688_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__a21oi_1
X_07399_ _02026_ _02028_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__xnor2_2
XFILLER_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09138_ sha256cu.iter_processing.w\[17\] _02639_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__nor2_1
XFILLER_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09069_ _03553_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__nand2_1
X_11100_ _04725_ _04721_ _04958_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__or3b_2
XFILLER_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12080_ sha256cu.data_in_padd\[20\] _05667_ _05892_ _05445_ VGND VGND VPWR VPWR _05893_
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11031_ sha256cu.data_in_padd\[5\] _01961_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__or2_1
XFILLER_134_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12982_ _02111_ _04917_ _05159_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__or3_2
X_11933_ _05751_ _05749_ _05433_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14721_ clknet_leaf_99_clk _01235_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11864_ _05684_ _05685_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__nor2_1
XFILLER_73_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14652_ clknet_leaf_122_clk _01166_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13603_ clknet_leaf_87_clk _00149_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10815_ _04701_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__clkbuf_4
X_11795_ sha256cu.iter_processing.w\[8\] _05430_ _05619_ _05335_ VGND VGND VPWR VPWR
+ _00906_ sky130_fd_sc_hd__o211a_1
X_14583_ clknet_leaf_122_clk _01097_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10746_ _01994_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13534_ clknet_leaf_103_clk _00084_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10677_ _04529_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__clkbuf_4
X_13465_ _06742_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12416_ _01912_ _05312_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__or2_2
XFILLER_127_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13396_ _06699_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12347_ _04743_ _06140_ _06142_ _01913_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__a211oi_1
XFILLER_142_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12278_ sha256cu.msg_scheduler.mreg_1\[15\] sha256cu.msg_scheduler.mreg_1\[4\] VGND
+ VGND VPWR VPWR _06082_ sky130_fd_sc_hd__xor2_1
XFILLER_107_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14017_ clknet_leaf_40_clk _00563_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11229_ _04907_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__buf_4
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14919_ clknet_leaf_2_clk _01433_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08440_ _02304_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__xnor2_2
XFILLER_64_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08371_ _02932_ _02935_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__nand2_1
XFILLER_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07322_ _01965_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__buf_4
XFILLER_31_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07253_ net257 _01908_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__and2b_1
X_07184_ _01792_ _01634_ _01653_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09825_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__clkbuf_2
XFILLER_86_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09756_ sha256cu.msg_scheduler.mreg_13\[3\] _04086_ _04094_ _04090_ VGND VGND VPWR
+ VPWR _00386_ sky130_fd_sc_hd__o211a_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06968_ _01586_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__clkbuf_4
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ sha256cu.msg_scheduler.mreg_14\[5\] _04045_ _04055_ _04050_ VGND VGND VPWR
+ VPWR _00356_ sky130_fd_sc_hd__o211a_1
X_08707_ _02051_ _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__xor2_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ sha256cu.m_out_digest.c_in\[18\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[18\]
+ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__o22a_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06899_ _01592_ _01577_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__nand2_2
XFILLER_15_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08569_ _03165_ _03167_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__xnor2_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ sha256cu.msg_scheduler.mreg_9\[4\] _04567_ _04578_ _04570_ VGND VGND VPWR
+ VPWR _00752_ sky130_fd_sc_hd__o211a_1
XFILLER_23_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11580_ _01937_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__inv_2
X_10531_ sha256cu.msg_scheduler.mreg_9\[7\] _04534_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__or2_1
XFILLER_22_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13250_ sha256cu.m_pad_pars.block_512\[52\]\[5\] _06617_ VGND VGND VPWR VPWR _06623_
+ sky130_fd_sc_hd__and2_1
X_10462_ sha256cu.msg_scheduler.mreg_7\[9\] _04487_ _04499_ _04490_ VGND VGND VPWR
+ VPWR _00693_ sky130_fd_sc_hd__o211a_1
XFILLER_108_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12201_ sha256cu.data_in_padd\[25\] _05667_ _06008_ _05445_ VGND VGND VPWR VPWR _06009_
+ sky130_fd_sc_hd__a211o_1
X_10393_ sha256cu.msg_scheduler.mreg_6\[11\] _04448_ _04460_ _04451_ VGND VGND VPWR
+ VPWR _00663_ sky130_fd_sc_hd__o211a_1
XFILLER_135_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13181_ sha256cu.m_pad_pars.block_512\[48\]\[5\] _06580_ VGND VGND VPWR VPWR _06586_
+ sky130_fd_sc_hd__and2_1
XFILLER_150_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12132_ sha256cu.msg_scheduler.mreg_9\[23\] sha256cu.msg_scheduler.mreg_0\[23\] VGND
+ VGND VPWR VPWR _05942_ sky130_fd_sc_hd__nand2_1
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12063_ _05874_ _05875_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__and2_1
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11014_ sha256cu.m_pad_pars.block_512\[3\]\[4\] _04765_ _04774_ sha256cu.m_pad_pars.block_512\[7\]\[4\]
+ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__a22o_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12965_ _01986_ _05303_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__or2_2
X_11916_ sha256cu.msg_scheduler.mreg_1\[21\] _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14704_ clknet_leaf_0_clk _01218_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_351 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12896_ _01912_ _05305_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__or2_2
XANTENNA_395 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ sha256cu.msg_scheduler.mreg_9\[11\] sha256cu.msg_scheduler.mreg_0\[11\] VGND
+ VGND VPWR VPWR _05669_ sky130_fd_sc_hd__nand2_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ clknet_leaf_8_clk _01149_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_362 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_384 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_373 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11778_ _05600_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__xor2_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14566_ clknet_leaf_116_clk _01080_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10729_ sha256cu.msg_scheduler.mreg_11\[28\] _04640_ VGND VGND VPWR VPWR _04652_
+ sky130_fd_sc_hd__or2_1
XFILLER_14_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13517_ sha256cu.temp_case sha256cu.iter_processing.padding_done _02000_ VGND VGND
+ VPWR VPWR _01473_ sky130_fd_sc_hd__o21a_1
X_14497_ clknet_leaf_104_clk _01011_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13448_ _06732_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13379_ _06690_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07940_ _02538_ _02540_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__or2b_1
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07871_ sha256cu.m_out_digest.g_in\[13\] sha256cu.m_out_digest.f_in\[13\] sha256cu.m_out_digest.e_in\[13\]
+ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__mux2_2
XFILLER_110_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09610_ _02109_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__clkbuf_4
X_06822_ net85 net88 net87 net91 VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__or4_1
XFILLER_56_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09541_ sha256cu.m_out_digest.h_in\[31\] sha256cu.m_out_digest.d_in\[31\] VGND VGND
+ VPWR VPWR _04012_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09472_ _03944_ _03945_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__and2_1
XFILLER_51_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08423_ _03024_ _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08354_ _02000_ _02958_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__nand2_1
X_07305_ _01939_ sha256cu.byte_rdy _01946_ _01948_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__o31a_1
X_08285_ sha256cu.m_out_digest.a_in\[14\] sha256cu.m_out_digest.a_in\[5\] VGND VGND
+ VPWR VPWR _02891_ sky130_fd_sc_hd__xnor2_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07236_ _01892_ _01893_ _01895_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07167_ _01836_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07098_ _01578_ _01653_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__nor2_1
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09808_ sha256cu.msg_scheduler.mreg_14\[26\] _04120_ VGND VGND VPWR VPWR _04124_
+ sky130_fd_sc_hd__or2_1
XFILLER_86_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09739_ sha256cu.msg_scheduler.mreg_14\[28\] _04073_ _04084_ _04077_ VGND VGND VPWR
+ VPWR _00379_ sky130_fd_sc_hd__o211a_1
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12750_ sha256cu.m_pad_pars.block_512\[23\]\[3\] _06353_ VGND VGND VPWR VPWR _06357_
+ sky130_fd_sc_hd__and2_1
X_11701_ _05517_ _05519_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__nand2_1
XFILLER_91_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ sha256cu.m_pad_pars.block_512\[19\]\[3\] _06316_ VGND VGND VPWR VPWR _06320_
+ sky130_fd_sc_hd__and2_1
XFILLER_42_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11632_ sha256cu.data_in_padd\[1\] _05448_ _05462_ _05463_ VGND VGND VPWR VPWR _05464_
+ sky130_fd_sc_hd__a211o_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ clknet_leaf_108_clk _00934_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_512_block\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14351_ clknet_leaf_7_clk _00865_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13302_ _06650_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
X_11563_ _04801_ _05275_ sha256cu.m_pad_pars.block_512\[40\]\[7\] VGND VGND VPWR VPWR
+ _05399_ sky130_fd_sc_hd__a21oi_1
X_10514_ _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__buf_2
X_14282_ clknet_leaf_24_clk _00828_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11494_ sha256cu.data_in_padd\[25\] _04840_ _05334_ _05335_ VGND VGND VPWR VPWR _00888_
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10445_ sha256cu.msg_scheduler.mreg_7\[1\] _04487_ _04489_ _04490_ VGND VGND VPWR
+ VPWR _00685_ sky130_fd_sc_hd__o211a_1
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13233_ sha256cu.m_pad_pars.block_512\[51\]\[5\] _06608_ VGND VGND VPWR VPWR _06614_
+ sky130_fd_sc_hd__and2_1
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13164_ sha256cu.m_pad_pars.block_512\[47\]\[5\] _06571_ VGND VGND VPWR VPWR _06577_
+ sky130_fd_sc_hd__and2_1
X_10376_ sha256cu.msg_scheduler.mreg_6\[3\] _04448_ _04450_ _04451_ VGND VGND VPWR
+ VPWR _00655_ sky130_fd_sc_hd__o211a_1
X_12115_ sha256cu.msg_scheduler.mreg_14\[9\] sha256cu.msg_scheduler.mreg_14\[7\] VGND
+ VGND VPWR VPWR _05926_ sky130_fd_sc_hd__xor2_1
XFILLER_97_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13095_ sha256cu.m_pad_pars.block_512\[43\]\[5\] _06534_ VGND VGND VPWR VPWR _06540_
+ sky130_fd_sc_hd__and2_1
XFILLER_2_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12046_ _05858_ _05859_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__and2b_1
XFILLER_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13997_ clknet_leaf_56_clk _00543_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12948_ _06270_ _04817_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__nand2_2
XFILLER_19_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12879_ _02111_ _04705_ _04809_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__or3_2
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14618_ clknet_leaf_121_clk _01132_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14549_ clknet_leaf_9_clk _01063_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_08070_ _02644_ _02647_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__o21a_1
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07021_ _01607_ _01608_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__nand2_4
XFILLER_127_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08972_ _03457_ _03461_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__and2_1
XFILLER_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07923_ _02503_ _02501_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__or2b_1
X_07854_ _02402_ _02471_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__nand2_1
XFILLER_69_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06805_ _01475_ _01476_ _01481_ _01502_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__or4_1
X_07785_ _02365_ _02404_ _02362_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__o21a_1
XFILLER_83_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09524_ sha256cu.K\[30\] _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__xnor2_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09455_ sha256cu.m_out_digest.h_in\[28\] sha256cu.m_out_digest.d_in\[28\] VGND VGND
+ VPWR VPWR _03929_ sky130_fd_sc_hd__nand2_1
XFILLER_24_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08406_ _03007_ _03008_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09386_ _03826_ _03842_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__and3_1
X_08337_ _02936_ _02941_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08268_ _02839_ _02843_ _02837_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__o21bai_1
XFILLER_153_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07219_ _01733_ _01659_ _01690_ _01603_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__o2bb2a_1
X_10230_ _04314_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__buf_2
XFILLER_118_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08199_ _02382_ sha256cu.m_out_digest.a_in\[3\] VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10161_ _04314_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__buf_2
XFILLER_133_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10092_ sha256cu.msg_scheduler.mreg_3\[10\] _04282_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__or2_1
XFILLER_120_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13920_ clknet_leaf_44_clk _00466_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13851_ clknet_leaf_21_clk _00397_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13782_ clknet_leaf_64_clk _00328_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12802_ _06384_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10994_ sha256cu.m_pad_pars.block_512\[35\]\[2\] _04818_ _04855_ _04858_ VGND VGND
+ VPWR VPWR _04859_ sky130_fd_sc_hd__a211o_1
X_12733_ _06347_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__clkbuf_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12664_ sha256cu.m_pad_pars.block_512\[18\]\[3\] _06307_ VGND VGND VPWR VPWR _06311_
+ sky130_fd_sc_hd__and2_1
X_14403_ clknet_leaf_76_clk _00917_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12595_ _06274_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_1
X_11615_ _05432_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11546_ sha256cu.m_pad_pars.block_512\[20\]\[6\] _05294_ _05314_ sha256cu.m_pad_pars.block_512\[0\]\[6\]
+ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__a221o_1
X_14334_ clknet_leaf_124_clk _00848_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.m_size\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14265_ clknet_leaf_20_clk _00811_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_13216_ sha256cu.m_pad_pars.block_512\[50\]\[5\] _06599_ VGND VGND VPWR VPWR _06605_
+ sky130_fd_sc_hd__and2_1
XFILLER_7_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11477_ _05319_ _05297_ _05278_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__and3b_2
X_10428_ sha256cu.msg_scheduler.mreg_6\[26\] _04474_ _04480_ _04477_ VGND VGND VPWR
+ VPWR _00678_ sky130_fd_sc_hd__o211a_1
X_14196_ clknet_leaf_29_clk _00742_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10359_ _04414_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__clkbuf_2
XFILLER_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13147_ sha256cu.m_pad_pars.block_512\[46\]\[5\] _06562_ VGND VGND VPWR VPWR _06568_
+ sky130_fd_sc_hd__and2_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13078_ sha256cu.m_pad_pars.block_512\[42\]\[5\] _06525_ VGND VGND VPWR VPWR _06531_
+ sky130_fd_sc_hd__and2_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12029_ _05841_ _05842_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__a21o_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07570_ sha256cu.m_out_digest.e_in\[16\] sha256cu.m_out_digest.e_in\[11\] VGND VGND
+ VPWR VPWR _02195_ sky130_fd_sc_hd__xnor2_2
XFILLER_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09240_ _03689_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__inv_2
XFILLER_22_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09171_ _03649_ _03653_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__and2_1
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08122_ _02233_ _02732_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__nand2_1
XFILLER_30_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08053_ _02654_ _02652_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__or2b_1
XFILLER_134_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07004_ _01606_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__buf_2
XFILLER_143_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08955_ _03416_ _03446_ _03414_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a21oi_2
Xinput108 hash[197] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput119 hash[206] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
X_07906_ _02520_ _02521_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08886_ _03378_ _03379_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__nand2_1
XFILLER_96_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07837_ _02451_ _02454_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__xnor2_2
X_07768_ _02345_ _02348_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__o21a_1
XFILLER_112_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09507_ _03944_ _03957_ _03977_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__and3_1
X_07699_ _02285_ _02287_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__nor2_1
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _03906_ _03911_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__and2_1
XFILLER_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09369_ _02931_ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__xor2_1
XFILLER_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12380_ _06159_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__clkbuf_1
X_11400_ _04787_ _04993_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__nor2_1
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_70 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_81 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ sha256cu.data_in_padd\[17\] _04741_ _04742_ _05180_ VGND VGND VPWR VPWR _00880_
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14050_ clknet_leaf_39_clk _00596_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11262_ _04726_ _04951_ _05111_ _05113_ _04976_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__a32o_1
XFILLER_4_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10213_ sha256cu.msg_scheduler.mreg_4\[30\] _04348_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__or2_1
X_11193_ sha256cu.m_pad_pars.block_512\[50\]\[3\] _05008_ _04972_ sha256cu.m_pad_pars.block_512\[38\]\[3\]
+ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__a221o_1
X_13001_ _06490_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10144_ sha256cu.msg_scheduler.mreg_4\[0\] _04308_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__or2_1
XFILLER_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10075_ sha256cu.msg_scheduler.mreg_3\[3\] _04268_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__or2_1
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14952_ clknet_leaf_89_clk _01466_ VGND VGND VPWR VPWR sha256cu.K\[25\] sky130_fd_sc_hd__dfxtp_1
X_14883_ clknet_leaf_99_clk _01397_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13903_ clknet_leaf_96_clk _00449_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.counter_iteration\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13834_ clknet_leaf_76_clk _00380_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[29\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13765_ clknet_leaf_81_clk _00311_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10977_ sha256cu.m_pad_pars.block_512\[63\]\[1\] _01920_ _04738_ _04833_ sha256cu.m_pad_pars.block_512\[55\]\[1\]
+ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__a32o_1
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13696_ clknet_leaf_68_clk _00242_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[19\]
+ sky130_fd_sc_hd__dfxtp_4
X_12716_ _06338_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_1
X_12647_ sha256cu.m_pad_pars.block_512\[17\]\[3\] _06298_ VGND VGND VPWR VPWR _06302_
+ sky130_fd_sc_hd__and2_1
XFILLER_31_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12578_ sha256cu.m_pad_pars.block_512\[13\]\[3\] _06261_ VGND VGND VPWR VPWR _06265_
+ sky130_fd_sc_hd__and2_1
XFILLER_7_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11529_ sha256cu.m_pad_pars.block_512\[32\]\[5\] _05306_ _05318_ sha256cu.m_pad_pars.block_512\[8\]\[5\]
+ _05366_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__a221o_1
X_14317_ clknet_leaf_95_clk _00010_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14248_ clknet_leaf_26_clk _00794_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_14179_ clknet_leaf_35_clk _00725_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ sha256cu.m_out_digest.e_in\[2\] _02040_ _03239_ _02068_ VGND VGND VPWR VPWR
+ _00225_ sky130_fd_sc_hd__a211o_1
XFILLER_39_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ sha256cu.m_out_digest.d_in\[15\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[15\]
+ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__o22a_1
X_07622_ _02208_ _02206_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__or2b_1
XFILLER_94_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07553_ _02140_ _02142_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__nor2_1
XFILLER_81_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07484_ _01911_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__clkbuf_8
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09223_ sha256cu.iter_processing.w\[20\] _02740_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__and2_1
XFILLER_22_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09154_ _03608_ _03638_ _03606_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__a21bo_1
X_08105_ sha256cu.m_out_digest.h_in\[19\] _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09085_ _03569_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__nand2_1
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08036_ sha256cu.m_out_digest.h_in\[16\] _02602_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__nand2_1
Xinput90 hash[180] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09987_ sha256cu.msg_scheduler.mreg_1\[29\] _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__or2_1
X_08938_ _03428_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__or2b_1
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08869_ _03362_ _03363_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10900_ sha256cu.m_pad_pars.add_out3\[3\] sha256cu.m_pad_pars.add_out3\[2\] VGND
+ VGND VPWR VPWR _04767_ sky130_fd_sc_hd__and2b_1
X_11880_ _05697_ _05699_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__or2_1
XFILLER_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10831_ sha256cu.m_pad_pars.m_size\[8\] _04706_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__or2_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10762_ sha256cu.msg_scheduler.mreg_11\[10\] _04659_ _04670_ _04662_ VGND VGND VPWR
+ VPWR _00822_ sky130_fd_sc_hd__o211a_1
X_13550_ clknet_leaf_75_clk _00096_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13481_ _06752_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__clkbuf_1
X_12501_ _01986_ _04933_ _05130_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__or3_2
XFILLER_139_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10693_ sha256cu.msg_scheduler.mreg_10\[12\] _04620_ _04631_ _04623_ VGND VGND VPWR
+ VPWR _00792_ sky130_fd_sc_hd__o211a_1
X_12432_ _06186_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12363_ sha256cu.m_pad_pars.block_512\[0\]\[6\] _06144_ VGND VGND VPWR VPWR _06151_
+ sky130_fd_sc_hd__and2_1
X_14102_ clknet_leaf_33_clk _00648_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12294_ sha256cu.msg_scheduler.mreg_9\[30\] sha256cu.msg_scheduler.mreg_0\[30\] VGND
+ VGND VPWR VPWR _06097_ sky130_fd_sc_hd__or2_1
X_11314_ _04912_ _05159_ _05152_ _05125_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__o211a_2
X_14033_ clknet_leaf_40_clk _00579_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11245_ sha256cu.m_pad_pars.block_512\[14\]\[7\] _05095_ _05096_ VGND VGND VPWR VPWR
+ _05097_ sky130_fd_sc_hd__o21a_1
XFILLER_5_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11176_ sha256cu.m_pad_pars.block_512\[26\]\[2\] _04964_ _05014_ sha256cu.m_pad_pars.block_512\[18\]\[2\]
+ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__a22o_1
XFILLER_68_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10127_ sha256cu.msg_scheduler.mreg_3\[25\] _04308_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__or2_1
XFILLER_121_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10058_ sha256cu.msg_scheduler.mreg_1\[27\] _04260_ _04269_ _04264_ VGND VGND VPWR
+ VPWR _00519_ sky130_fd_sc_hd__o211a_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14935_ clknet_leaf_88_clk _01449_ VGND VGND VPWR VPWR sha256cu.K\[8\] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14866_ clknet_leaf_1_clk _01380_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13817_ clknet_leaf_48_clk _00363_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_14797_ clknet_leaf_11_clk _01311_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13748_ clknet_leaf_61_clk _00294_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13679_ clknet_leaf_72_clk _00225_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09910_ _04177_ _04184_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__nor2_1
XFILLER_113_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09841_ sha256cu.msg_scheduler.mreg_13\[8\] _04134_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__or2_1
XFILLER_86_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ sha256cu.msg_scheduler.mreg_13\[10\] _04099_ _04102_ _04103_ VGND VGND VPWR
+ VPWR _00393_ sky130_fd_sc_hd__o211a_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _01669_ _01671_ _01620_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__mux2_1
X_08723_ sha256cu.iter_processing.w\[2\] _02075_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__or2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ sha256cu.m_out_digest.d_in\[1\] _03185_ _03186_ sha256cu.m_out_digest.c_in\[1\]
+ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__o22a_1
X_08585_ sha256cu.m_out_digest.b_in\[7\] _02370_ _02110_ sha256cu.m_out_digest.a_in\[7\]
+ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__o22a_1
X_07605_ sha256cu.m_out_digest.e_in\[17\] sha256cu.m_out_digest.e_in\[12\] VGND VGND
+ VPWR VPWR _02229_ sky130_fd_sc_hd__xnor2_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07536_ sha256cu.m_out_digest.a_in\[17\] VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07467_ _02092_ _02094_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__xnor2_1
X_09206_ _03657_ _03669_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__and3_1
XFILLER_136_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07398_ _02027_ sha256cu.m_out_digest.a_in\[2\] VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__xnor2_1
X_09137_ _03620_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__xnor2_1
X_09068_ _03502_ _03554_ _03555_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__o21bai_1
XFILLER_118_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08019_ _02612_ _02614_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__or2b_1
XFILLER_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11030_ _04887_ _04889_ _04890_ _04891_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__or4_2
XFILLER_2_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12981_ _06479_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__clkbuf_1
X_11932_ _05704_ _05707_ _05725_ _05724_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__a31o_1
X_14720_ clknet_leaf_99_clk _01234_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11863_ _05658_ _05662_ _05683_ _05432_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__a31o_1
XFILLER_60_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14651_ clknet_leaf_123_clk _01165_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13602_ clknet_leaf_86_clk _00148_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10814_ sha256cu.m_pad_pars.temp_chk VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__clkbuf_4
X_11794_ sha256cu.data_in_padd\[8\] _05433_ _05616_ _05618_ _04046_ VGND VGND VPWR
+ VPWR _05619_ sky130_fd_sc_hd__a221o_1
X_14582_ clknet_leaf_113_clk _01096_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10745_ sha256cu.msg_scheduler.mreg_12\[3\] _04653_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__or2_1
XFILLER_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13533_ clknet_leaf_107_clk _00083_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10676_ sha256cu.msg_scheduler.mreg_11\[5\] _04614_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__or2_1
X_13464_ _06730_ _06741_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__and2_1
XFILLER_145_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12415_ _06177_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__clkbuf_1
X_13395_ sha256cu.m_pad_pars.block_512\[61\]\[2\] _06693_ VGND VGND VPWR VPWR _06699_
+ sky130_fd_sc_hd__and2_1
XFILLER_9_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12346_ sha256cu.byte_rdy _01914_ _04777_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__and3_1
XFILLER_153_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12277_ _06079_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__nand2_1
X_14016_ clknet_leaf_40_clk _00562_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11228_ sha256cu.data_in_padd\[14\] _04840_ _05078_ _05080_ _05040_ VGND VGND VPWR
+ VPWR _00877_ sky130_fd_sc_hd__o221a_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11159_ sha256cu.m_pad_pars.block_512\[6\]\[0\] _04957_ _04965_ _05017_ VGND VGND
+ VPWR VPWR _05018_ sky130_fd_sc_hd__a211o_1
XFILLER_83_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14918_ clknet_leaf_117_clk _01432_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14849_ clknet_leaf_99_clk _01363_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ _02968_ _02973_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07321_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__buf_6
XFILLER_16_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07252_ state\[1\] sha256cu.hashing_done _01560_ net258 VGND VGND VPWR VPWR _01908_
+ sky130_fd_sc_hd__a31o_1
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07183_ _01657_ _01687_ _01849_ _01633_ _01621_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__a221o_1
XFILLER_129_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09824_ _01566_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__buf_4
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09755_ sha256cu.msg_scheduler.mreg_14\[3\] _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__or2_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06967_ _01607_ _01642_ _01653_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__a31o_1
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09686_ sha256cu.iter_processing.w\[5\] _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__or2_1
X_08706_ _03205_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__nand2_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06898_ _01573_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__clkinv_2
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ sha256cu.m_out_digest.c_in\[17\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[17\]
+ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__o22a_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08568_ sha256cu.m_out_digest.a_in\[21\] _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__xnor2_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07519_ _02115_ _02116_ _02144_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__a21oi_2
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08499_ _03097_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10530_ sha256cu.msg_scheduler.mreg_8\[6\] _04526_ _04538_ _04530_ VGND VGND VPWR
+ VPWR _00722_ sky130_fd_sc_hd__o211a_1
XFILLER_129_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10461_ sha256cu.msg_scheduler.mreg_8\[9\] _04494_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__or2_1
XFILLER_109_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12200_ _06005_ _06006_ _06007_ _05442_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__o211a_1
X_10392_ sha256cu.msg_scheduler.mreg_7\[11\] _04455_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__or2_1
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13180_ _06585_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__clkbuf_1
X_12131_ sha256cu.msg_scheduler.mreg_9\[23\] sha256cu.msg_scheduler.mreg_0\[23\] VGND
+ VGND VPWR VPWR _05941_ sky130_fd_sc_hd__or2_1
XFILLER_108_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12062_ _05872_ _05873_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__nand2_1
XFILLER_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11013_ sha256cu.m_pad_pars.block_512\[27\]\[4\] _04757_ _04804_ sha256cu.m_pad_pars.block_512\[43\]\[4\]
+ _04875_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__a221o_1
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12964_ _06470_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11915_ sha256cu.msg_scheduler.mreg_1\[17\] sha256cu.msg_scheduler.mreg_1\[0\] VGND
+ VGND VPWR VPWR _05734_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14703_ clknet_leaf_0_clk _01217_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_352 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_330 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12895_ _06433_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_385 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ sha256cu.msg_scheduler.mreg_9\[11\] sha256cu.msg_scheduler.mreg_0\[11\] VGND
+ VGND VPWR VPWR _05668_ sky130_fd_sc_hd__or2_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ clknet_leaf_16_clk _01148_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_374 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_363 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_396 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11777_ sha256cu.msg_scheduler.mreg_1\[26\] _05601_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__xnor2_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14565_ clknet_leaf_98_clk _01079_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10728_ sha256cu.msg_scheduler.mreg_10\[27\] _04646_ _04651_ _04649_ VGND VGND VPWR
+ VPWR _00807_ sky130_fd_sc_hd__o211a_1
X_13516_ _06774_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14496_ clknet_leaf_105_clk _01010_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10659_ sha256cu.msg_scheduler.mreg_9\[29\] _04607_ _04612_ _04610_ VGND VGND VPWR
+ VPWR _00777_ sky130_fd_sc_hd__o211a_1
X_13447_ _06730_ _06731_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__and2_1
XFILLER_142_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13378_ sha256cu.m_pad_pars.block_512\[60\]\[2\] _06682_ VGND VGND VPWR VPWR _06690_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12329_ sha256cu.iter_processing.w\[31\] _04044_ _06129_ _06130_ _05040_ VGND VGND
+ VPWR VPWR _00929_ sky130_fd_sc_hd__o221a_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07870_ sha256cu.m_out_digest.b_in\[13\] _02027_ _02486_ VGND VGND VPWR VPWR _02487_
+ sky130_fd_sc_hd__o21ai_1
X_06821_ net76 net80 net79 net82 VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__or4_1
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09540_ sha256cu.K\[30\] _03995_ _03994_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09471_ _03904_ _03912_ _03943_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__or3_1
XFILLER_64_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08422_ _02981_ _02985_ _03023_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__or3b_1
XFILLER_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08353_ sha256cu.m_out_digest.a_in\[25\] _02629_ _02923_ _02957_ VGND VGND VPWR VPWR
+ _02958_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07304_ _01939_ _01947_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__nand2_1
X_08284_ _02856_ _02861_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__nand2_1
XFILLER_20_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07235_ _01652_ _01761_ _01894_ _01570_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__o31a_1
XFILLER_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07166_ _01833_ _01835_ _01570_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__mux2_1
X_07097_ _01646_ _01634_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__nor2_1
XFILLER_59_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07999_ _02574_ _02576_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__and2_1
XFILLER_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09807_ sha256cu.msg_scheduler.mreg_13\[25\] _04112_ _04123_ _04117_ VGND VGND VPWR
+ VPWR _00408_ sky130_fd_sc_hd__o211a_1
XFILLER_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09738_ sha256cu.iter_processing.w\[28\] _04080_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__or2_1
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__buf_6
X_11700_ _05526_ _05527_ _05528_ _05335_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__o211a_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12680_ _06319_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__clkbuf_1
X_11631_ _04053_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__buf_2
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14350_ clknet_leaf_9_clk _00864_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11562_ _01935_ _05297_ _05394_ _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__a31o_1
X_10513_ _01972_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__buf_2
X_13301_ sha256cu.m_pad_pars.block_512\[55\]\[5\] _06644_ VGND VGND VPWR VPWR _06650_
+ sky130_fd_sc_hd__and2_1
XFILLER_109_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14281_ clknet_leaf_25_clk _00827_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11493_ _01994_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10444_ _04396_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__buf_2
XFILLER_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13232_ _06613_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10375_ _04396_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__buf_2
XFILLER_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ _06576_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12114_ _05923_ _05924_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__and2_1
XFILLER_124_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13094_ _06539_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__clkbuf_1
X_12045_ _05828_ _05833_ _05857_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__a21o_1
XFILLER_2_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13996_ clknet_leaf_57_clk _00542_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12947_ _01966_ _05121_ _06461_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12878_ _06424_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_160 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11829_ sha256cu.msg_scheduler.mreg_14\[27\] sha256cu.msg_scheduler.mreg_14\[20\]
+ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__xnor2_1
XANTENNA_171 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14617_ clknet_leaf_121_clk _01131_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14548_ clknet_leaf_6_clk _01062_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14479_ clknet_leaf_6_clk _00993_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_07020_ _01701_ _01704_ _01596_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__o21ai_4
XFILLER_114_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08971_ _03457_ _03461_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__nor2_1
X_07922_ _02518_ _02537_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07853_ _02401_ _02435_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__and2b_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06804_ _01486_ _01491_ _01496_ _01501_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__or4_1
XFILLER_68_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07784_ _02334_ _02361_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__nor2_1
XFILLER_37_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09523_ _03993_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__nor2_1
XFILLER_37_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09454_ _03890_ _03919_ _03920_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__o21ba_1
XFILLER_24_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08405_ sha256cu.m_out_digest.g_in\[27\] sha256cu.m_out_digest.f_in\[27\] sha256cu.m_out_digest.e_in\[27\]
+ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09385_ _03860_ _03861_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08336_ sha256cu.iter_processing.w\[25\] _02940_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__xor2_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08267_ _02871_ _02873_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__xor2_2
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08198_ sha256cu.K\[22\] VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__inv_2
X_07218_ _01684_ _01820_ _01799_ _01585_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__a211o_1
XFILLER_146_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07149_ _01603_ _01610_ _01706_ _01820_ _01620_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__a311o_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10160_ sha256cu.msg_scheduler.mreg_3\[7\] _04315_ _04327_ _04318_ VGND VGND VPWR
+ VPWR _00563_ sky130_fd_sc_hd__o211a_1
XFILLER_133_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10091_ _04166_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__buf_2
XFILLER_126_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13850_ clknet_leaf_17_clk _00396_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13781_ clknet_leaf_65_clk _00327_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_90_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12801_ sha256cu.m_pad_pars.block_512\[26\]\[3\] _06380_ VGND VGND VPWR VPWR _06384_
+ sky130_fd_sc_hd__and2_1
XFILLER_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10993_ sha256cu.m_pad_pars.block_512\[43\]\[2\] _04804_ _04828_ sha256cu.m_pad_pars.block_512\[23\]\[2\]
+ _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__a221o_1
X_12732_ sha256cu.m_pad_pars.block_512\[22\]\[3\] _06343_ VGND VGND VPWR VPWR _06347_
+ sky130_fd_sc_hd__and2_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14402_ clknet_leaf_75_clk _00916_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_12663_ _06310_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__clkbuf_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ sha256cu.iter_processing.w\[0\] _05430_ _05446_ _05335_ VGND VGND VPWR VPWR
+ _00898_ sky130_fd_sc_hd__o211a_1
X_12594_ sha256cu.m_pad_pars.block_512\[14\]\[2\] _06271_ VGND VGND VPWR VPWR _06274_
+ sky130_fd_sc_hd__and2_1
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11545_ sha256cu.m_pad_pars.block_512\[28\]\[6\] _05296_ _05381_ _01920_ VGND VGND
+ VPWR VPWR _05382_ sky130_fd_sc_hd__a22o_1
X_14333_ clknet_leaf_2_clk _00847_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.m_size\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14264_ clknet_leaf_27_clk _00810_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11476_ _05275_ _05316_ _04801_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__o21a_1
X_10427_ sha256cu.msg_scheduler.mreg_7\[26\] _04468_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__or2_1
X_13215_ _06604_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__clkbuf_1
X_14195_ clknet_leaf_29_clk _00741_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10358_ sha256cu.msg_scheduler.mreg_5\[28\] _04434_ _04440_ _04437_ VGND VGND VPWR
+ VPWR _00648_ sky130_fd_sc_hd__o211a_1
XFILLER_97_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13146_ _06567_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__clkbuf_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _04281_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__clkbuf_2
XFILLER_112_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13077_ _06530_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12028_ sha256cu.data_in_padd\[18\] _05447_ _04692_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__a21o_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13979_ clknet_leaf_54_clk _00525_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09170_ _03649_ _03653_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__nor2_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08121_ _02037_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_122_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_30_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08052_ _02662_ _02663_ _02664_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07003_ _00453_ _01589_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__nor2_2
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput109 hash[198] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
X_08954_ _03394_ _03395_ _03412_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__a21o_1
XFILLER_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07905_ sha256cu.m_out_digest.g_in\[14\] sha256cu.m_out_digest.f_in\[14\] sha256cu.m_out_digest.e_in\[14\]
+ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__mux2_1
X_08885_ sha256cu.iter_processing.w\[8\] _02296_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__or2_1
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07836_ sha256cu.m_out_digest.h_in\[12\] _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__xnor2_2
XFILLER_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07767_ sha256cu.m_out_digest.h_in\[9\] _02347_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__nand2_1
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09506_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__inv_2
XFILLER_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07698_ sha256cu.K\[8\] _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__xnor2_2
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ _03906_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__nor2_1
XFILLER_40_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ _03843_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__nand2_1
XFILLER_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09299_ _03777_ _03778_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_113_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_16
X_08319_ sha256cu.K\[25\] VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__inv_2
XANTENNA_71 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _05172_ _05174_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__or3_1
XANTENNA_60 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11261_ _04801_ _04974_ _05112_ sha256cu.m_pad_pars.block_512\[46\]\[7\] VGND VGND
+ VPWR VPWR _05113_ sky130_fd_sc_hd__a22o_1
X_10212_ sha256cu.msg_scheduler.mreg_3\[29\] _04354_ _04356_ _04357_ VGND VGND VPWR
+ VPWR _00585_ sky130_fd_sc_hd__o211a_1
XFILLER_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11192_ sha256cu.m_pad_pars.block_512\[34\]\[3\] _04996_ _04981_ sha256cu.m_pad_pars.block_512\[54\]\[3\]
+ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__a22o_1
X_13000_ sha256cu.m_pad_pars.block_512\[38\]\[0\] _06489_ VGND VGND VPWR VPWR _06490_
+ sky130_fd_sc_hd__and2_1
X_10143_ sha256cu.msg_scheduler.mreg_2\[31\] _04315_ _04317_ _04318_ VGND VGND VPWR
+ VPWR _00555_ sky130_fd_sc_hd__o211a_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10074_ sha256cu.msg_scheduler.mreg_2\[2\] _04274_ _04278_ _04277_ VGND VGND VPWR
+ VPWR _00526_ sky130_fd_sc_hd__o211a_1
XFILLER_102_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14951_ clknet_leaf_90_clk _01465_ VGND VGND VPWR VPWR sha256cu.K\[24\] sky130_fd_sc_hd__dfxtp_2
XFILLER_101_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14882_ clknet_leaf_101_clk _01396_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13902_ clknet_leaf_95_clk _00448_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.counter_iteration\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13833_ clknet_leaf_110_clk _00379_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[28\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13764_ clknet_leaf_85_clk _00310_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10976_ sha256cu.m_pad_pars.block_512\[3\]\[1\] _04765_ _04841_ _01970_ VGND VGND
+ VPWR VPWR _04842_ sky130_fd_sc_hd__a211o_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13695_ clknet_leaf_68_clk _00241_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[18\]
+ sky130_fd_sc_hd__dfxtp_4
X_12715_ sha256cu.m_pad_pars.block_512\[21\]\[3\] _06334_ VGND VGND VPWR VPWR _06338_
+ sky130_fd_sc_hd__and2_1
XFILLER_31_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12646_ _06301_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_104_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_16
X_12577_ _06264_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14316_ clknet_leaf_92_clk _00009_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__dfxtp_1
X_11528_ sha256cu.m_pad_pars.block_512\[24\]\[5\] _05279_ _05304_ sha256cu.m_pad_pars.block_512\[36\]\[5\]
+ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__a22o_1
X_14247_ clknet_leaf_26_clk _00793_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11459_ _04794_ _05154_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__nor2_1
X_14178_ clknet_leaf_35_clk _00724_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13129_ _06558_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__clkbuf_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08670_ sha256cu.m_out_digest.d_in\[14\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[14\]
+ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__o22a_1
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07621_ _02221_ _02244_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__xnor2_2
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07552_ sha256cu.K\[4\] _02177_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07483_ _02070_ _02106_ _02107_ _02110_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__a2bb2o_1
X_09222_ sha256cu.iter_processing.w\[20\] _02740_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__nor2_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09153_ _03612_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__inv_2
XFILLER_147_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08104_ sha256cu.m_out_digest.a_in\[21\] _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09084_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__inv_2
X_08035_ _02644_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__xnor2_1
Xinput91 hash[181] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
Xinput80 hash[171] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09986_ _04133_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__clkbuf_2
XFILLER_89_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08937_ _03426_ _03427_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nand2_1
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08868_ _03336_ _03339_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__nand2_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07819_ _02435_ _02437_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__xnor2_2
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08799_ _03294_ _03295_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10830_ sha256cu.m_pad_pars.add_512_block\[4\] _04700_ _04712_ _04709_ VGND VGND
+ VPWR VPWR _00848_ sky130_fd_sc_hd__o211a_1
X_10761_ sha256cu.msg_scheduler.mreg_12\[10\] _04666_ VGND VGND VPWR VPWR _04670_
+ sky130_fd_sc_hd__or2_1
X_10692_ sha256cu.msg_scheduler.mreg_11\[12\] _04627_ VGND VGND VPWR VPWR _04631_
+ sky130_fd_sc_hd__or2_1
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12500_ _06222_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
X_13480_ _06730_ _06751_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__and2_1
X_12431_ sha256cu.m_pad_pars.block_512\[4\]\[7\] _05411_ _01983_ VGND VGND VPWR VPWR
+ _06186_ sky130_fd_sc_hd__mux2_1
XFILLER_148_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12362_ _06150_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14101_ clknet_leaf_33_clk _00647_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12293_ sha256cu.iter_processing.w\[29\] _05894_ _06096_ _01974_ VGND VGND VPWR VPWR
+ _00927_ sky130_fd_sc_hd__o211a_1
XFILLER_4_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11313_ sha256cu.m_pad_pars.block_512\[61\]\[0\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[0\]
+ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__a22o_1
X_14032_ clknet_leaf_40_clk _00578_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11244_ _04786_ _04973_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__nand2_1
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11175_ sha256cu.m_pad_pars.block_512\[6\]\[2\] _04957_ _04989_ sha256cu.m_pad_pars.block_512\[14\]\[2\]
+ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__a221o_1
X_10126_ _04281_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10057_ sha256cu.msg_scheduler.mreg_2\[27\] _04268_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__or2_1
XFILLER_0_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14934_ clknet_leaf_89_clk _01448_ VGND VGND VPWR VPWR sha256cu.K\[7\] sky130_fd_sc_hd__dfxtp_4
XFILLER_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14865_ clknet_leaf_1_clk _01379_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13816_ clknet_leaf_48_clk _00362_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_14796_ clknet_leaf_14_clk _01310_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13747_ clknet_leaf_60_clk _00293_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10959_ _04823_ _04825_ _04736_ _04764_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__and4bb_4
XFILLER_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13678_ clknet_leaf_71_clk _00224_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12629_ _06292_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09840_ sha256cu.msg_scheduler.mreg_12\[7\] _04140_ _04142_ _04130_ VGND VGND VPWR
+ VPWR _00422_ sky130_fd_sc_hd__o211a_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09771_ _01973_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__buf_2
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _01670_ _01661_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__xnor2_1
X_08722_ sha256cu.iter_processing.w\[2\] _02075_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__nand2_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _02109_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__buf_4
XFILLER_27_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07604_ sha256cu.iter_processing.w\[6\] _02227_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__xnor2_2
X_08584_ sha256cu.m_out_digest.b_in\[6\] _03031_ _02114_ sha256cu.m_out_digest.a_in\[6\]
+ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__a22o_1
XFILLER_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07535_ sha256cu.m_out_digest.a_in\[26\] VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__buf_4
XFILLER_53_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07466_ _02049_ _02059_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09205_ _03686_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07397_ sha256cu.m_out_digest.a_in\[13\] VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09136_ _02599_ _03585_ _03586_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__a21boi_1
XFILLER_136_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09067_ _03496_ _03526_ _03525_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08018_ _02128_ _02220_ _02628_ _02631_ _02258_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__a221o_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09969_ sha256cu.msg_scheduler.mreg_0\[21\] _04208_ _04218_ _04211_ VGND VGND VPWR
+ VPWR _00481_ sky130_fd_sc_hd__o211a_1
XFILLER_134_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12980_ sha256cu.m_pad_pars.block_512\[36\]\[7\] _05401_ _06442_ VGND VGND VPWR VPWR
+ _06479_ sky130_fd_sc_hd__mux2_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _05704_ _05707_ _05725_ _05749_ _05724_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__a311o_4
XFILLER_27_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11862_ _05658_ _05662_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__a21oi_1
X_14650_ clknet_leaf_123_clk _01164_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13601_ clknet_leaf_85_clk _00147_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10813_ _04698_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__nand2_2
X_14581_ clknet_leaf_4_clk _01095_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11793_ _05447_ _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__nor2_1
X_13532_ clknet_leaf_107_clk _00082_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out1\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10744_ sha256cu.msg_scheduler.mreg_11\[2\] _04659_ _04660_ _04649_ VGND VGND VPWR
+ VPWR _00814_ sky130_fd_sc_hd__o211a_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10675_ sha256cu.msg_scheduler.mreg_10\[4\] _04620_ _04621_ _04610_ VGND VGND VPWR
+ VPWR _00784_ sky130_fd_sc_hd__o211a_1
X_13463_ sha256cu.K\[12\] _06714_ _06719_ _00039_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__a22o_1
X_12414_ sha256cu.m_pad_pars.block_512\[3\]\[7\] _04935_ _01983_ VGND VGND VPWR VPWR
+ _06177_ sky130_fd_sc_hd__mux2_1
X_13394_ _06698_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12345_ _06141_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12276_ sha256cu.msg_scheduler.mreg_9\[29\] sha256cu.msg_scheduler.mreg_0\[29\] VGND
+ VGND VPWR VPWR _06080_ sky130_fd_sc_hd__or2_1
X_14015_ clknet_leaf_56_clk _00561_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11227_ sha256cu.m_pad_pars.block_512\[18\]\[6\] _05014_ _05079_ _01970_ VGND VGND
+ VPWR VPWR _05080_ sky130_fd_sc_hd__a211o_1
XFILLER_150_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11158_ sha256cu.m_pad_pars.block_512\[38\]\[0\] _04972_ _04986_ _05003_ _05016_
+ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__a2111o_1
X_10109_ sha256cu.msg_scheduler.mreg_2\[17\] _04288_ _04298_ _04291_ VGND VGND VPWR
+ VPWR _00541_ sky130_fd_sc_hd__o211a_1
XFILLER_110_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11089_ _04756_ _04764_ _04943_ _04948_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__a31o_1
XFILLER_64_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14917_ clknet_leaf_99_clk _01431_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14848_ clknet_leaf_99_clk _01362_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07320_ _01564_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__clkbuf_4
X_14779_ clknet_leaf_125_clk _01293_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_07251_ _01907_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07182_ _00452_ _01640_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nand2_1
XFILLER_8_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09823_ sha256cu.msg_scheduler.mreg_12\[0\] _04126_ _04132_ _04130_ VGND VGND VPWR
+ VPWR _00415_ sky130_fd_sc_hd__o211a_1
XFILLER_100_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09754_ _04053_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__clkbuf_2
X_06966_ _01654_ _01590_ _01634_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__and3_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08705_ sha256cu.m_out_digest.h_in\[1\] sha256cu.m_out_digest.d_in\[1\] VGND VGND
+ VPWR VPWR _03206_ sky130_fd_sc_hd__or2_1
X_09685_ _04053_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__clkbuf_2
XFILLER_73_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06897_ _01586_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__nor2_2
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08636_ _02369_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__buf_4
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ sha256cu.K\[31\] sha256cu.m_out_digest.h_in\[31\] VGND VGND VPWR VPWR _03166_
+ sky130_fd_sc_hd__xor2_1
X_07518_ _02115_ _02116_ _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__nand3_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08498_ sha256cu.iter_processing.w\[28\] _03053_ _03098_ VGND VGND VPWR VPWR _03099_
+ sky130_fd_sc_hd__a21oi_1
X_07449_ _02073_ _02074_ _02075_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__a21o_1
XFILLER_136_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10460_ sha256cu.msg_scheduler.mreg_7\[8\] _04487_ _04498_ _04490_ VGND VGND VPWR
+ VPWR _00692_ sky130_fd_sc_hd__o211a_1
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09119_ _03576_ _03577_ _03604_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__a21bo_1
X_10391_ sha256cu.msg_scheduler.mreg_6\[10\] _04448_ _04459_ _04451_ VGND VGND VPWR
+ VPWR _00662_ sky130_fd_sc_hd__o211a_1
XFILLER_124_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12130_ sha256cu.iter_processing.w\[22\] _05894_ _05940_ _05866_ VGND VGND VPWR VPWR
+ _00920_ sky130_fd_sc_hd__o211a_1
XFILLER_2_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12061_ _05872_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__or2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11012_ sha256cu.m_pad_pars.block_512\[51\]\[4\] _04826_ _04822_ sha256cu.m_pad_pars.block_512\[47\]\[4\]
+ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__a221o_1
XFILLER_104_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12963_ sha256cu.m_pad_pars.block_512\[35\]\[7\] _04920_ _06442_ VGND VGND VPWR VPWR
+ _06470_ sky130_fd_sc_hd__mux2_1
XFILLER_18_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _05731_ _05732_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_84_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
X_14702_ clknet_leaf_111_clk _01216_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_320 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_331 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14633_ clknet_leaf_16_clk _01147_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_342 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12894_ sha256cu.m_pad_pars.block_512\[31\]\[7\] _04911_ _06351_ VGND VGND VPWR VPWR
+ _06433_ sky130_fd_sc_hd__mux2_1
XANTENNA_353 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11845_ _05447_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__clkbuf_4
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_364 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_386 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_397 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11776_ sha256cu.msg_scheduler.mreg_1\[15\] sha256cu.msg_scheduler.mreg_1\[11\] VGND
+ VGND VPWR VPWR _05601_ sky130_fd_sc_hd__xnor2_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ clknet_leaf_96_clk _01078_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10727_ sha256cu.msg_scheduler.mreg_11\[27\] _04640_ VGND VGND VPWR VPWR _04651_
+ sky130_fd_sc_hd__or2_1
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14495_ clknet_leaf_104_clk _01009_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13515_ _01975_ _06773_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__and2_1
XFILLER_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13446_ sha256cu.K\[5\] _06714_ _06719_ _00063_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__a22o_1
X_10658_ sha256cu.msg_scheduler.mreg_10\[29\] _04601_ VGND VGND VPWR VPWR _04612_
+ sky130_fd_sc_hd__or2_1
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10589_ sha256cu.msg_scheduler.mreg_8\[31\] _04567_ _04572_ _04570_ VGND VGND VPWR
+ VPWR _00747_ sky130_fd_sc_hd__o211a_1
XFILLER_115_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13377_ _06689_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12328_ sha256cu.data_in_padd\[31\] _05448_ _05463_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__a21o_1
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12259_ _06062_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__or2_2
XFILLER_69_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06820_ net81 net84 net83 net86 VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__or4_1
XFILLER_49_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
X_09470_ _03904_ _03912_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08421_ _02981_ _02985_ _03023_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__o21ba_1
XFILLER_24_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08352_ _02955_ _02956_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__xnor2_1
X_07303_ sha256cu.byte_stop _01916_ sha256cu.byte_rdy VGND VGND VPWR VPWR _01947_
+ sky130_fd_sc_hd__a21o_1
X_08283_ _02855_ _02852_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__or2b_1
XFILLER_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07234_ _01607_ _01580_ _01646_ _00452_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__o211a_1
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07165_ _01703_ _01831_ _01834_ _01617_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__o22a_1
XFILLER_105_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07096_ _01618_ _01771_ _01772_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__a22o_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07998_ _02592_ _02611_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__xnor2_1
X_09806_ sha256cu.msg_scheduler.mreg_14\[25\] _04120_ VGND VGND VPWR VPWR _04123_
+ sky130_fd_sc_hd__or2_1
XFILLER_28_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09737_ sha256cu.msg_scheduler.mreg_14\[27\] _04073_ _04083_ _04077_ VGND VGND VPWR
+ VPWR _00378_ sky130_fd_sc_hd__o211a_1
X_06949_ _01588_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_66_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09668_ sha256cu.msg_scheduler.counter_iteration\[5\] sha256cu.msg_scheduler.counter_iteration\[4\]
+ _01565_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__or3_1
X_08619_ sha256cu.m_out_digest.c_in\[3\] _03179_ _03178_ sha256cu.m_out_digest.b_in\[3\]
+ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__a22o_1
X_09599_ sha256cu.m_out_digest.g_in\[3\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[3\]
+ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__o22a_1
XFILLER_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _05460_ _05461_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__nor2_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11561_ _05277_ _05293_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__and3_1
X_10512_ sha256cu.msg_scheduler.mreg_8\[31\] _04520_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__or2_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13300_ _06649_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
X_14280_ clknet_leaf_25_clk _00826_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11492_ sha256cu.m_pad_pars.block_512\[0\]\[1\] _05314_ _05333_ _01971_ VGND VGND
+ VPWR VPWR _05334_ sky130_fd_sc_hd__a211o_1
XFILLER_136_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10443_ sha256cu.msg_scheduler.mreg_8\[1\] _04481_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__or2_1
X_13231_ sha256cu.m_pad_pars.block_512\[51\]\[4\] _06608_ VGND VGND VPWR VPWR _06613_
+ sky130_fd_sc_hd__and2_1
X_10374_ sha256cu.msg_scheduler.mreg_7\[3\] _04441_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__or2_1
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13162_ sha256cu.m_pad_pars.block_512\[47\]\[4\] _06571_ VGND VGND VPWR VPWR _06576_
+ sky130_fd_sc_hd__and2_1
XFILLER_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12113_ _05921_ _05922_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__nand2_1
XFILLER_151_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13093_ sha256cu.m_pad_pars.block_512\[43\]\[4\] _06534_ VGND VGND VPWR VPWR _06539_
+ sky130_fd_sc_hd__and2_1
XFILLER_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12044_ _05828_ _05833_ _05857_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__and3_1
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13995_ clknet_leaf_57_clk _00541_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_57_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_46_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12946_ _03288_ sha256cu.m_pad_pars.block_512\[34\]\[7\] VGND VGND VPWR VPWR _06461_
+ sky130_fd_sc_hd__nor2_1
XFILLER_45_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_150 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ sha256cu.m_pad_pars.block_512\[30\]\[7\] _05102_ _06351_ VGND VGND VPWR VPWR
+ _06424_ sky130_fd_sc_hd__mux2_1
XANTENNA_161 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11828_ _05649_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__and2_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14616_ clknet_leaf_120_clk _01130_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ clknet_leaf_5_clk _01061_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11759_ _05582_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__xor2_1
X_14478_ clknet_leaf_113_clk _00992_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13429_ _06718_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08970_ sha256cu.K\[11\] _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__xor2_1
XFILLER_88_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07921_ _02534_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07852_ _02467_ _02469_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__xor2_1
XFILLER_96_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput1 hash[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_06803_ _01497_ _01498_ _01499_ _01500_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__or4_1
XFILLER_68_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07783_ _02402_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_48_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
X_09522_ sha256cu.iter_processing.w\[30\] _03126_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__and2_1
XFILLER_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09453_ _03839_ _03895_ _03925_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__o31a_1
XFILLER_52_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08404_ sha256cu.m_out_digest.b_in\[27\] sha256cu.m_out_digest.a_in\[27\] _03006_
+ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__o21ai_1
XFILLER_52_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09384_ sha256cu.K\[24\] _03823_ _03822_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__a21o_1
XFILLER_61_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08335_ _02938_ _02939_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08266_ _02806_ _02835_ _02872_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__o21ai_2
X_08197_ _02792_ _02794_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__or2b_1
X_07217_ _01595_ _01604_ _01751_ _01618_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__o31ai_1
XFILLER_146_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07148_ _01743_ _01639_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__and2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07079_ _01632_ _01617_ _01721_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__or3_1
X_10090_ sha256cu.msg_scheduler.mreg_2\[9\] _04274_ _04287_ _04277_ VGND VGND VPWR
+ VPWR _00533_ sky130_fd_sc_hd__o211a_1
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12800_ _06383_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__clkbuf_1
X_13780_ clknet_leaf_61_clk _00326_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_83_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10992_ sha256cu.m_pad_pars.block_512\[27\]\[2\] _04757_ _04790_ sha256cu.m_pad_pars.block_512\[11\]\[2\]
+ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__a221o_1
XFILLER_16_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12731_ _06346_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__clkbuf_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12662_ sha256cu.m_pad_pars.block_512\[18\]\[2\] _06307_ VGND VGND VPWR VPWR _06310_
+ sky130_fd_sc_hd__and2_1
XFILLER_70_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11613_ sha256cu.data_in_padd\[0\] _05433_ _05443_ _05444_ _05445_ VGND VGND VPWR
+ VPWR _05446_ sky130_fd_sc_hd__a221o_1
X_14401_ clknet_leaf_75_clk _00915_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12593_ _06273_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11544_ sha256cu.m_pad_pars.block_512\[60\]\[6\] _01998_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[6\]
+ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__a22o_1
X_14332_ clknet_leaf_2_clk _00846_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.m_size\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14263_ clknet_leaf_20_clk _00809_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11475_ _05315_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nor2_4
X_10426_ sha256cu.msg_scheduler.mreg_6\[25\] _04474_ _04479_ _04477_ VGND VGND VPWR
+ VPWR _00677_ sky130_fd_sc_hd__o211a_1
X_13214_ sha256cu.m_pad_pars.block_512\[50\]\[4\] _06599_ VGND VGND VPWR VPWR _06604_
+ sky130_fd_sc_hd__and2_1
XFILLER_136_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14194_ clknet_leaf_29_clk _00740_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10357_ sha256cu.msg_scheduler.mreg_6\[28\] _04428_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__or2_1
X_13145_ sha256cu.m_pad_pars.block_512\[46\]\[4\] _06562_ VGND VGND VPWR VPWR _06567_
+ sky130_fd_sc_hd__and2_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ sha256cu.msg_scheduler.mreg_4\[30\] _04393_ _04400_ _04397_ VGND VGND VPWR
+ VPWR _00618_ sky130_fd_sc_hd__o211a_1
XFILLER_112_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13076_ sha256cu.m_pad_pars.block_512\[42\]\[4\] _06525_ VGND VGND VPWR VPWR _06530_
+ sky130_fd_sc_hd__and2_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12027_ _05840_ _05818_ _05820_ _05433_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__a31oi_1
XFILLER_93_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13978_ clknet_leaf_42_clk _00524_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12929_ sha256cu.m_pad_pars.block_512\[33\]\[7\] _05267_ _06442_ VGND VGND VPWR VPWR
+ _06452_ sky130_fd_sc_hd__mux2_1
XFILLER_33_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08120_ _02728_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__xor2_1
X_08051_ _02162_ _02440_ _01966_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__o21ai_1
X_07002_ _01654_ _01687_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__nor2_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08953_ _03391_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__nor2_1
XFILLER_103_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07904_ sha256cu.m_out_digest.b_in\[14\] sha256cu.m_out_digest.a_in\[14\] _02519_
+ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08884_ sha256cu.iter_processing.w\[8\] _02296_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__nand2_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07835_ sha256cu.m_out_digest.a_in\[25\] _02452_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__xnor2_2
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07766_ _02381_ _02385_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09505_ _03944_ _03957_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a21o_1
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07697_ _02316_ _02318_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__xnor2_2
X_09436_ sha256cu.K\[27\] _03910_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__xnor2_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09367_ sha256cu.m_out_digest.h_in\[25\] sha256cu.m_out_digest.d_in\[25\] VGND VGND
+ VPWR VPWR _03844_ sky130_fd_sc_hd__nand2_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_50 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08318_ _02065_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__clkbuf_4
X_09298_ _03744_ _03756_ _03776_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__nand3_1
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_72 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08249_ _02852_ _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__xnor2_1
XANTENNA_61 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_94 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11260_ _04801_ _04973_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__nand2_1
X_10211_ _04263_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__buf_2
X_11191_ _05041_ _05044_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__or3_1
X_10142_ _04263_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__clkbuf_4
X_10073_ sha256cu.msg_scheduler.mreg_3\[2\] _04268_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__or2_1
XFILLER_95_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14950_ clknet_leaf_89_clk _01464_ VGND VGND VPWR VPWR sha256cu.K\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14881_ clknet_leaf_99_clk _01395_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13901_ clknet_leaf_95_clk _00447_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.counter_iteration\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13832_ clknet_leaf_76_clk _00378_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[27\]
+ sky130_fd_sc_hd__dfxtp_2
X_13763_ clknet_leaf_84_clk _00309_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10975_ sha256cu.m_pad_pars.block_512\[7\]\[1\] _04774_ _04781_ sha256cu.m_pad_pars.block_512\[15\]\[1\]
+ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__a22o_1
XFILLER_43_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ _06337_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_1
X_13694_ clknet_leaf_67_clk _00240_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[17\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12645_ sha256cu.m_pad_pars.block_512\[17\]\[2\] _06298_ VGND VGND VPWR VPWR _06301_
+ sky130_fd_sc_hd__and2_1
X_12576_ sha256cu.m_pad_pars.block_512\[13\]\[2\] _06261_ VGND VGND VPWR VPWR _06264_
+ sky130_fd_sc_hd__and2_1
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11527_ sha256cu.data_in_padd\[28\] _01980_ _01987_ _05365_ VGND VGND VPWR VPWR _00891_
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14315_ clknet_leaf_91_clk _00008_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14246_ clknet_leaf_27_clk _00792_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11458_ sha256cu.m_pad_pars.block_512\[20\]\[0\] _05294_ _05296_ sha256cu.m_pad_pars.block_512\[28\]\[0\]
+ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__a221o_1
X_10409_ sha256cu.msg_scheduler.mreg_7\[18\] _04468_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__or2_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14177_ clknet_leaf_35_clk _00723_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11389_ _04704_ _05154_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__or2_1
XFILLER_98_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13128_ sha256cu.m_pad_pars.block_512\[45\]\[4\] _06553_ VGND VGND VPWR VPWR _06558_
+ sky130_fd_sc_hd__and2_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13059_ sha256cu.m_pad_pars.block_512\[41\]\[4\] _06516_ VGND VGND VPWR VPWR _06521_
+ sky130_fd_sc_hd__and2_1
XFILLER_78_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07620_ _02241_ _02243_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__xnor2_2
X_07551_ _02174_ _02176_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__xor2_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07482_ _02109_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__buf_4
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09221_ _03701_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__or2_1
XFILLER_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09152_ _03635_ _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__and2b_1
XFILLER_147_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08103_ sha256cu.m_out_digest.a_in\[9\] sha256cu.m_out_digest.a_in\[0\] VGND VGND
+ VPWR VPWR _02714_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09083_ sha256cu.iter_processing.w\[15\] _02561_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__and2_1
Xinput70 hash[162] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
Xinput81 hash[172] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
XFILLER_147_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08034_ sha256cu.m_out_digest.h_in\[17\] _02646_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__xnor2_1
Xinput92 hash[182] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
X_09985_ sha256cu.msg_scheduler.mreg_0\[28\] _04221_ _04227_ _04224_ VGND VGND VPWR
+ VPWR _00488_ sky130_fd_sc_hd__o211a_1
XFILLER_107_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08936_ _03426_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__nor2_1
XFILLER_103_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08867_ _03360_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__or2b_1
XFILLER_111_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07818_ _02401_ _02406_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__o21ba_1
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ _02159_ _03265_ _03266_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__a21boi_1
XFILLER_84_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07749_ _02017_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__clkbuf_4
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10760_ sha256cu.msg_scheduler.mreg_11\[9\] _04659_ _04669_ _04662_ VGND VGND VPWR
+ VPWR _00821_ sky130_fd_sc_hd__o211a_1
XFILLER_80_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10691_ sha256cu.msg_scheduler.mreg_10\[11\] _04620_ _04630_ _04623_ VGND VGND VPWR
+ VPWR _00791_ sky130_fd_sc_hd__o211a_1
X_09419_ _03834_ _03865_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__or2b_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12430_ _06185_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14100_ clknet_leaf_37_clk _00646_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12361_ sha256cu.m_pad_pars.block_512\[0\]\[5\] _06144_ VGND VGND VPWR VPWR _06150_
+ sky130_fd_sc_hd__and2_1
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12292_ _05442_ _06093_ _06094_ _06095_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__a31o_1
X_11312_ _05139_ _05149_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__and2_2
X_14031_ clknet_leaf_40_clk _00577_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11243_ _04702_ _04780_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nor2_1
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11174_ sha256cu.m_pad_pars.block_512\[2\]\[2\] _04999_ _05030_ _01921_ VGND VGND
+ VPWR VPWR _05031_ sky130_fd_sc_hd__a22o_1
X_10125_ sha256cu.msg_scheduler.mreg_2\[24\] _04301_ _04307_ _04304_ VGND VGND VPWR
+ VPWR _00548_ sky130_fd_sc_hd__o211a_1
X_10056_ _04133_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__clkbuf_2
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14933_ clknet_leaf_89_clk _01447_ VGND VGND VPWR VPWR sha256cu.K\[6\] sky130_fd_sc_hd__dfxtp_4
XFILLER_75_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14864_ clknet_leaf_1_clk _01378_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13815_ clknet_leaf_48_clk _00361_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14795_ clknet_leaf_13_clk _01309_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13746_ clknet_leaf_60_clk _00292_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10958_ _04761_ _04824_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__nor2_2
X_13677_ clknet_leaf_72_clk _00223_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_92_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10889_ _04735_ sha256cu.m_pad_pars.add_out3\[4\] VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__and2_2
X_12628_ sha256cu.m_pad_pars.block_512\[16\]\[2\] _06289_ VGND VGND VPWR VPWR _06292_
+ sky130_fd_sc_hd__and2_1
XFILLER_12_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12559_ sha256cu.m_pad_pars.block_512\[12\]\[2\] _06252_ VGND VGND VPWR VPWR _06255_
+ sky130_fd_sc_hd__and2_1
X_14229_ clknet_leaf_27_clk _00775_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[27\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_125_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ sha256cu.msg_scheduler.mreg_14\[10\] _04093_ VGND VGND VPWR VPWR _04102_
+ sky130_fd_sc_hd__or2_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ _01632_ _01649_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__nor2_1
X_08721_ _03211_ _03214_ _03212_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ sha256cu.m_out_digest.d_in\[0\] _03184_ _03182_ sha256cu.m_out_digest.c_in\[0\]
+ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__a22o_1
XFILLER_66_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07603_ _02225_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__and2b_1
X_08583_ sha256cu.m_out_digest.b_in\[5\] _03031_ _02114_ sha256cu.m_out_digest.a_in\[5\]
+ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__a22o_1
XFILLER_82_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07534_ _02159_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__inv_2
X_07465_ _02056_ _02058_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__nor2_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09204_ sha256cu.K\[18\] _03652_ _03651_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__a21o_1
XFILLER_10_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07396_ sha256cu.m_out_digest.a_in\[22\] VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__buf_4
X_09135_ _02643_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__xor2_1
X_09066_ _03498_ _03527_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__or2b_1
XFILLER_135_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08017_ _02629_ _02630_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__nor2_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09968_ sha256cu.msg_scheduler.mreg_1\[21\] _04215_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__or2_1
XFILLER_103_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08919_ _03410_ _03411_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11930_ _05747_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__nand2_1
XFILLER_73_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09899_ _01564_ sha256cu.iter_processing.padding_done VGND VGND VPWR VPWR _04177_
+ sky130_fd_sc_hd__nand2_2
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11861_ _05681_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__or2b_1
X_11792_ _05593_ _05594_ _05597_ _05615_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__and4_1
X_13600_ clknet_leaf_84_clk _00146_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_14580_ clknet_leaf_4_clk _01094_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10812_ sha256cu.byte_rdy _01945_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__nor2_8
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10743_ sha256cu.msg_scheduler.mreg_12\[2\] _04653_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__or2_1
X_13531_ clknet_leaf_107_clk _00081_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out1\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_41_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10674_ sha256cu.msg_scheduler.mreg_11\[4\] _04614_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__or2_1
X_13462_ sha256cu.K\[11\] _06726_ _06727_ _06740_ _06737_ VGND VGND VPWR VPWR _01452_
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12413_ _06176_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__clkbuf_1
X_13393_ sha256cu.m_pad_pars.block_512\[61\]\[1\] _06693_ VGND VGND VPWR VPWR _06698_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12344_ _01973_ _06139_ _06140_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__and3_1
XFILLER_153_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14014_ clknet_leaf_41_clk _00560_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12275_ sha256cu.msg_scheduler.mreg_9\[29\] sha256cu.msg_scheduler.mreg_0\[29\] VGND
+ VGND VPWR VPWR _06079_ sky130_fd_sc_hd__nand2_1
XFILLER_5_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11226_ sha256cu.m_pad_pars.block_512\[42\]\[6\] _05001_ _05013_ sha256cu.m_pad_pars.block_512\[22\]\[6\]
+ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__a22o_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11157_ sha256cu.m_pad_pars.block_512\[50\]\[0\] _05008_ _05009_ sha256cu.m_pad_pars.block_512\[30\]\[0\]
+ _05015_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__a221o_1
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10108_ sha256cu.msg_scheduler.mreg_3\[17\] _04295_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__or2_1
XFILLER_110_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11088_ _04755_ _04756_ _04945_ _04946_ _04947_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__a32o_1
X_10039_ sha256cu.msg_scheduler.mreg_2\[20\] _04254_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__or2_1
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14916_ clknet_leaf_100_clk _01430_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14847_ clknet_leaf_98_clk _01361_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14778_ clknet_leaf_121_clk _01292_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13729_ clknet_leaf_83_clk _00275_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07250_ sha256cu.byte_stop _01906_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__and2_1
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07181_ _01687_ _01719_ _01702_ _01703_ _01585_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__a221o_1
XFILLER_118_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09822_ sha256cu.msg_scheduler.mreg_13\[0\] _04120_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__or2_1
XFILLER_140_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09753_ sha256cu.msg_scheduler.mreg_13\[2\] _04086_ _04092_ _04090_ VGND VGND VPWR
+ VPWR _00385_ sky130_fd_sc_hd__o211a_1
XFILLER_59_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08704_ sha256cu.m_out_digest.h_in\[1\] sha256cu.m_out_digest.d_in\[1\] VGND VGND
+ VPWR VPWR _03205_ sky130_fd_sc_hd__nand2_1
X_06965_ _01608_ _01648_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__or2_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09684_ _01566_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06896_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__buf_4
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ sha256cu.m_out_digest.c_in\[16\] _03184_ _03182_ sha256cu.m_out_digest.b_in\[16\]
+ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__a22o_1
XFILLER_82_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08566_ sha256cu.m_out_digest.b_in\[31\] sha256cu.m_out_digest.a_in\[31\] _03164_
+ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__o21a_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07517_ sha256cu.K\[3\] _02143_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__xnor2_1
X_08497_ _03051_ _03052_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__and2b_1
X_07448_ _02073_ _02074_ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__and3_1
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07379_ Hash_Digest _02010_ _02012_ _02000_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__o211a_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09118_ _03575_ _03574_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__or2b_1
X_10390_ sha256cu.msg_scheduler.mreg_7\[10\] _04455_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__or2_1
XFILLER_135_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09049_ _02492_ _03509_ _03508_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12060_ _05845_ _05849_ _05846_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__a21boi_1
XFILLER_2_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11011_ sha256cu.m_pad_pars.block_512\[31\]\[4\] _04811_ _04872_ _04738_ _04873_
+ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__a221o_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12962_ _06469_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__clkbuf_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ sha256cu.msg_scheduler.mreg_9\[14\] sha256cu.msg_scheduler.mreg_0\[14\] VGND
+ VGND VPWR VPWR _05732_ sky130_fd_sc_hd__nand2_1
XANTENNA_310 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14701_ clknet_leaf_22_clk _01215_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12893_ _06432_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__clkbuf_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11844_ _04043_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14632_ clknet_leaf_12_clk _01146_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_343 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_332 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_376 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_365 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_354 net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_398 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11775_ _05598_ _05599_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__nand2_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_387 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14563_ clknet_leaf_96_clk _01077_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ sha256cu.msg_scheduler.mreg_10\[26\] _04646_ _04650_ _04649_ VGND VGND VPWR
+ VPWR _00806_ sky130_fd_sc_hd__o211a_1
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14494_ clknet_leaf_123_clk _01008_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13514_ sha256cu.K\[31\] _06713_ _06718_ _00060_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__a22o_1
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10657_ sha256cu.msg_scheduler.mreg_9\[28\] _04607_ _04611_ _04610_ VGND VGND VPWR
+ VPWR _00776_ sky130_fd_sc_hd__o211a_1
XFILLER_9_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13445_ _01972_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__buf_2
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10588_ sha256cu.msg_scheduler.mreg_9\[31\] _04561_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__or2_1
X_13376_ sha256cu.m_pad_pars.block_512\[60\]\[1\] _06682_ VGND VGND VPWR VPWR _06689_
+ sky130_fd_sc_hd__and2_1
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12327_ _06127_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__nor2_1
XFILLER_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12258_ _06033_ _06037_ _06034_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__a21boi_1
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11209_ _05024_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__and2_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12189_ _05994_ _05995_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__nand2_1
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08420_ _02996_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08351_ _02885_ _02920_ _02918_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__o21ba_1
XFILLER_60_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07302_ _01942_ _01944_ _01945_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__a21oi_1
X_08282_ sha256cu.K\[24\] VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__inv_2
X_07233_ _01739_ _01809_ _00456_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07164_ _01580_ _01602_ _01830_ _01747_ _01608_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__o32a_1
X_07095_ _01657_ _01646_ _01696_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__or3_1
XFILLER_132_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07997_ _02608_ _02610_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__xnor2_1
X_09805_ sha256cu.msg_scheduler.mreg_13\[24\] _04112_ _04122_ _04117_ VGND VGND VPWR
+ VPWR _00407_ sky130_fd_sc_hd__o211a_1
XFILLER_75_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09736_ sha256cu.iter_processing.w\[27\] _04080_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__or2_1
X_06948_ _01578_ _01637_ _01612_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__and3_1
X_09667_ sha256cu.m_out_digest.h_in\[31\] _04041_ _02113_ sha256cu.m_out_digest.g_in\[31\]
+ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__a22o_1
X_08618_ sha256cu.m_out_digest.c_in\[2\] _03179_ _03178_ sha256cu.m_out_digest.b_in\[2\]
+ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a22o_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06879_ sha256cu.iter_processing.rst _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nand2_8
XFILLER_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09598_ sha256cu.m_out_digest.g_in\[2\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[2\]
+ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__a22o_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08549_ sha256cu.K\[30\] _03139_ _03138_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__a21oi_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11560_ _04747_ _04815_ _05395_ sha256cu.m_pad_pars.block_512\[20\]\[7\] VGND VGND
+ VPWR VPWR _05396_ sky130_fd_sc_hd__o22a_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10511_ sha256cu.msg_scheduler.mreg_7\[30\] _04526_ _04527_ _04516_ VGND VGND VPWR
+ VPWR _00714_ sky130_fd_sc_hd__o211a_1
X_11491_ _05327_ _05328_ _05330_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__or4_1
X_13230_ _06612_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10442_ sha256cu.msg_scheduler.mreg_7\[0\] _04487_ _04488_ _04477_ VGND VGND VPWR
+ VPWR _00684_ sky130_fd_sc_hd__o211a_1
XFILLER_109_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10373_ sha256cu.msg_scheduler.mreg_6\[2\] _04448_ _04449_ _04437_ VGND VGND VPWR
+ VPWR _00654_ sky130_fd_sc_hd__o211a_1
XFILLER_123_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13161_ _06575_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12112_ _05921_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__or2_1
X_13092_ _06538_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12043_ _05854_ _05856_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13994_ clknet_leaf_58_clk _00540_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12945_ _06460_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_151 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _06423_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_140 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _05647_ _05648_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__nand2_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14615_ clknet_leaf_123_clk _01129_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11758_ _05583_ _05560_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__nand2_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ clknet_leaf_3_clk _01060_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_195 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10709_ sha256cu.msg_scheduler.mreg_11\[19\] _04640_ VGND VGND VPWR VPWR _04641_
+ sky130_fd_sc_hd__or2_1
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11689_ sha256cu.msg_scheduler.mreg_14\[21\] sha256cu.msg_scheduler.mreg_14\[14\]
+ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__xnor2_1
X_14477_ clknet_leaf_8_clk _00991_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13428_ sha256cu.counter_iteration\[6\] _06717_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__nor2_4
XFILLER_127_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13359_ sha256cu.m_pad_pars.block_512\[59\]\[1\] _06671_ VGND VGND VPWR VPWR _06680_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07920_ _02490_ _02500_ _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__o21ba_1
X_07851_ sha256cu.K\[11\] _02433_ _02468_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__a21o_1
XFILLER_111_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07782_ _02323_ _02362_ _02363_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__and3b_1
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06802_ net239 net242 net241 net244 VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__or4_1
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 hash[100] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09521_ sha256cu.iter_processing.w\[30\] _03126_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__nor2_1
XFILLER_37_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _03896_ _03925_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__or2_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08403_ sha256cu.m_out_digest.b_in\[27\] sha256cu.m_out_digest.a_in\[27\] sha256cu.m_out_digest.c_in\[27\]
+ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__a21o_1
XFILLER_52_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09383_ _03858_ _03859_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__xnor2_1
X_08334_ sha256cu.m_out_digest.g_in\[25\] sha256cu.m_out_digest.f_in\[25\] sha256cu.m_out_digest.e_in\[25\]
+ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__mux2_1
XFILLER_138_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08265_ _02832_ _02834_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__or2b_1
XFILLER_20_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08196_ _02332_ _02803_ _02804_ _02000_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__o211a_1
XFILLER_20_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07216_ _01679_ _01875_ _01876_ _01878_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__o22a_1
X_07147_ _01690_ _01750_ _01682_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__and3_1
XFILLER_133_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07078_ _01722_ _01757_ _01644_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__a21o_1
XFILLER_87_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09719_ _04044_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__buf_2
X_10991_ sha256cu.m_pad_pars.block_512\[63\]\[2\] _01920_ _04738_ _04833_ sha256cu.m_pad_pars.block_512\[55\]\[2\]
+ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__a32o_1
X_12730_ sha256cu.m_pad_pars.block_512\[22\]\[2\] _06343_ VGND VGND VPWR VPWR _06346_
+ sky130_fd_sc_hd__and2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12661_ _06309_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__clkbuf_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14400_ clknet_leaf_75_clk _00914_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_11612_ _04053_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__clkbuf_4
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12592_ sha256cu.m_pad_pars.block_512\[14\]\[1\] _06271_ VGND VGND VPWR VPWR _06273_
+ sky130_fd_sc_hd__and2_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11543_ sha256cu.m_pad_pars.block_512\[16\]\[6\] _05285_ _05288_ sha256cu.m_pad_pars.block_512\[48\]\[6\]
+ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__a22o_1
X_14331_ clknet_leaf_114_clk _00845_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.m_size\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14262_ clknet_leaf_27_clk _00808_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11474_ _05275_ _05316_ _04786_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__o21a_1
XFILLER_143_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10425_ sha256cu.msg_scheduler.mreg_7\[25\] _04468_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__or2_1
X_14193_ clknet_leaf_29_clk _00739_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_13213_ _06603_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13144_ _06566_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10356_ sha256cu.msg_scheduler.mreg_5\[27\] _04434_ _04439_ _04437_ VGND VGND VPWR
+ VPWR _00647_ sky130_fd_sc_hd__o211a_1
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ sha256cu.msg_scheduler.mreg_5\[30\] _04387_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__or2_1
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13075_ _06529_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _05818_ _05820_ _05840_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__a21o_1
XFILLER_120_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13977_ clknet_leaf_42_clk _00523_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[31\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12928_ _06451_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__clkbuf_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _06414_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14529_ clknet_leaf_106_clk _01043_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08050_ _02619_ _02630_ _02661_ _02515_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__o31a_1
XFILLER_134_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07001_ _01640_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08952_ _03389_ _03415_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__nand2_1
XFILLER_130_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08883_ sha256cu.K\[8\] VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__inv_2
X_07903_ sha256cu.m_out_digest.b_in\[14\] sha256cu.m_out_digest.a_in\[14\] sha256cu.m_out_digest.c_in\[14\]
+ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__a21o_1
XFILLER_97_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07834_ sha256cu.m_out_digest.a_in\[14\] sha256cu.m_out_digest.a_in\[2\] VGND VGND
+ VPWR VPWR _02452_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07765_ sha256cu.m_out_digest.h_in\[10\] _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07696_ _02261_ _02284_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__a21bo_1
X_09504_ _03975_ _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09435_ _03908_ _03909_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__nor2_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ sha256cu.m_out_digest.h_in\[25\] sha256cu.m_out_digest.d_in\[25\] VGND VGND
+ VPWR VPWR _03843_ sky130_fd_sc_hd__or2_1
XANTENNA_40 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ _03744_ _03756_ _03776_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__a21o_1
X_08317_ _02113_ _02921_ _02922_ _02332_ _02083_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__a32o_1
XANTENNA_73 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _02853_ _02811_ _02854_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__a21oi_1
XANTENNA_62 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_95 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ sha256cu.msg_scheduler.mreg_4\[29\] _04348_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__or2_1
X_08179_ _02782_ _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11190_ sha256cu.m_pad_pars.block_512\[10\]\[3\] _04963_ _05001_ sha256cu.m_pad_pars.block_512\[42\]\[3\]
+ _05045_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__a221o_1
X_10141_ sha256cu.msg_scheduler.mreg_3\[31\] _04308_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__or2_1
XFILLER_121_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10072_ sha256cu.msg_scheduler.mreg_2\[1\] _04274_ _04276_ _04277_ VGND VGND VPWR
+ VPWR _00525_ sky130_fd_sc_hd__o211a_1
X_13900_ clknet_leaf_18_clk _00446_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14880_ clknet_leaf_99_clk _01394_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13831_ clknet_leaf_76_clk _00377_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[26\]
+ sky130_fd_sc_hd__dfxtp_2
X_13762_ clknet_leaf_84_clk _00308_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10974_ _01963_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__buf_4
XFILLER_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12713_ sha256cu.m_pad_pars.block_512\[21\]\[2\] _06334_ VGND VGND VPWR VPWR _06337_
+ sky130_fd_sc_hd__and2_1
X_13693_ clknet_leaf_68_clk _00239_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[16\]
+ sky130_fd_sc_hd__dfxtp_4
X_12644_ _06300_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__clkbuf_1
X_12575_ _06263_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11526_ _05357_ _05359_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__or3_2
X_14314_ clknet_leaf_92_clk _00007_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14245_ clknet_leaf_27_clk _00791_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11457_ sha256cu.m_pad_pars.block_512\[44\]\[0\] _05298_ _05299_ sha256cu.m_pad_pars.block_512\[12\]\[0\]
+ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__a22o_1
X_10408_ sha256cu.msg_scheduler.mreg_6\[17\] _04461_ _04469_ _04464_ VGND VGND VPWR
+ VPWR _00669_ sky130_fd_sc_hd__o211a_1
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14176_ clknet_leaf_35_clk _00722_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11388_ _04917_ _05129_ _05231_ sha256cu.m_pad_pars.block_512\[41\]\[7\] VGND VGND
+ VPWR VPWR _05232_ sky130_fd_sc_hd__o22a_1
X_10339_ sha256cu.msg_scheduler.mreg_6\[20\] _04428_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__or2_1
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _06557_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _06520_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12009_ sha256cu.msg_scheduler.mreg_1\[21\] sha256cu.msg_scheduler.mreg_1\[4\] VGND
+ VGND VPWR VPWR _05824_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07550_ _02117_ _02139_ _02175_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07481_ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__buf_2
X_09220_ _03699_ _03700_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__and2_1
XFILLER_34_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09151_ _03615_ _03616_ _03634_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__a21o_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09082_ sha256cu.iter_processing.w\[15\] _02561_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__or2_1
X_08102_ _02712_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__inv_2
XFILLER_147_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08033_ _02304_ _02645_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__xnor2_2
Xinput82 hash[173] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xinput60 hash[153] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
Xinput71 hash[163] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xinput93 hash[183] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_143_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09984_ sha256cu.msg_scheduler.mreg_1\[28\] _04215_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__or2_1
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08935_ _02344_ _03396_ _03397_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__a21boi_1
XFILLER_85_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08866_ _03329_ _03341_ _03359_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__a21o_1
X_07817_ _02398_ _02400_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__nor2_1
X_08797_ _02196_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07748_ sha256cu.m_out_digest.a_in\[9\] _02040_ _02368_ _02068_ VGND VGND VPWR VPWR
+ _00104_ sky130_fd_sc_hd__a211o_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07679_ sha256cu.m_out_digest.e_in\[14\] sha256cu.m_out_digest.e_in\[1\] VGND VGND
+ VPWR VPWR _02301_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10690_ sha256cu.msg_scheduler.mreg_11\[11\] _04627_ VGND VGND VPWR VPWR _04630_
+ sky130_fd_sc_hd__or2_1
X_09418_ _03840_ _03869_ _03893_ _03863_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__a211o_1
XFILLER_13_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09349_ _03791_ _03799_ _03825_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__or3_1
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12360_ _06149_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11311_ _01977_ _05149_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__and2_2
X_12291_ sha256cu.data_in_padd\[29\] _05447_ _04053_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__a21o_1
XFILLER_153_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14030_ clknet_leaf_40_clk _00576_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11242_ _04726_ _04958_ _05083_ _05089_ _05093_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__a311o_1
X_11173_ sha256cu.m_pad_pars.block_512\[62\]\[2\] _04984_ _04982_ sha256cu.m_pad_pars.block_512\[58\]\[2\]
+ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__a22o_1
X_10124_ sha256cu.msg_scheduler.mreg_3\[24\] _04295_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__or2_1
XFILLER_121_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10055_ sha256cu.msg_scheduler.mreg_1\[26\] _04260_ _04267_ _04264_ VGND VGND VPWR
+ VPWR _00518_ sky130_fd_sc_hd__o211a_1
XFILLER_76_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14932_ clknet_leaf_95_clk _01446_ VGND VGND VPWR VPWR sha256cu.K\[5\] sky130_fd_sc_hd__dfxtp_4
XFILLER_76_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14863_ clknet_leaf_1_clk _01377_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13814_ clknet_leaf_47_clk _00360_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_75_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14794_ clknet_leaf_12_clk _01308_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13745_ clknet_leaf_66_clk _00291_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10957_ _01956_ _01914_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__nand2_4
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13676_ clknet_leaf_71_clk _00222_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10888_ sha256cu.m_pad_pars.add_out3\[2\] sha256cu.m_pad_pars.add_out3\[3\] VGND
+ VGND VPWR VPWR _04755_ sky130_fd_sc_hd__and2b_1
X_12627_ _06291_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__clkbuf_1
X_12558_ _06254_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__clkbuf_1
X_12489_ sha256cu.m_pad_pars.block_512\[8\]\[2\] _06214_ VGND VGND VPWR VPWR _06217_
+ sky130_fd_sc_hd__and2_1
X_11509_ sha256cu.m_pad_pars.block_512\[12\]\[3\] _05299_ _05304_ sha256cu.m_pad_pars.block_512\[36\]\[3\]
+ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__a221o_1
X_14228_ clknet_leaf_26_clk _00774_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[26\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_153_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14159_ clknet_leaf_31_clk _00705_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _01646_ _01666_ _01668_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08720_ _03202_ _03216_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__nand2_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ sha256cu.m_out_digest.c_in\[31\] _03184_ _03182_ sha256cu.m_out_digest.b_in\[31\]
+ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__a22o_1
XFILLER_82_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07602_ _02222_ _02223_ _02224_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__a21o_1
XFILLER_94_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08582_ sha256cu.m_out_digest.b_in\[4\] _03031_ _02114_ sha256cu.m_out_digest.a_in\[4\]
+ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__a22o_1
X_07533_ sha256cu.m_out_digest.e_in\[29\] _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__xnor2_2
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07464_ _02079_ _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__xor2_1
X_09203_ _03684_ _03685_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__nor2_1
X_07395_ _02024_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__inv_2
X_09134_ _03617_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__nand2_1
XFILLER_50_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09065_ _03551_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__and2_1
X_08016_ _02621_ _02627_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__nor2_2
XFILLER_144_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09967_ sha256cu.msg_scheduler.mreg_0\[20\] _04208_ _04217_ _04211_ VGND VGND VPWR
+ VPWR _00480_ sky130_fd_sc_hd__o211a_1
X_08918_ _03377_ _03380_ _03378_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__o21ai_1
XFILLER_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ sha256cu.msg_scheduler.counter_iteration\[0\] sha256cu.msg_scheduler.temp_case
+ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__and2_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _03321_ _03327_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__nor2_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11860_ _05649_ _05654_ _05680_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__a21o_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11791_ _05593_ _05594_ _05597_ _05615_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__a31o_1
X_10811_ _01956_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__clkbuf_4
XFILLER_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10742_ _04580_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__clkbuf_4
X_13530_ clknet_leaf_108_clk _00080_ VGND VGND VPWR VPWR sha256cu.byte_rdy sky130_fd_sc_hd__dfxtp_2
XFILLER_53_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10673_ _04580_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__buf_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13461_ _04188_ _00038_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__and2b_1
XFILLER_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12412_ sha256cu.m_pad_pars.block_512\[3\]\[6\] _06169_ VGND VGND VPWR VPWR _06176_
+ sky130_fd_sc_hd__and2_1
X_13392_ _06697_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ sha256cu.m_pad_pars.add_512_block\[4\] _06136_ VGND VGND VPWR VPWR _06140_
+ sky130_fd_sc_hd__nand2_1
X_12274_ sha256cu.iter_processing.w\[28\] _05894_ _06078_ _05866_ VGND VGND VPWR VPWR
+ _00926_ sky130_fd_sc_hd__o211a_1
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14013_ clknet_leaf_41_clk _00559_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11225_ sha256cu.m_pad_pars.block_512\[10\]\[6\] _04963_ _04996_ sha256cu.m_pad_pars.block_512\[34\]\[6\]
+ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__a221o_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11156_ sha256cu.m_pad_pars.block_512\[22\]\[0\] _05013_ _05014_ sha256cu.m_pad_pars.block_512\[18\]\[0\]
+ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__a22o_1
X_10107_ sha256cu.msg_scheduler.mreg_2\[16\] _04288_ _04297_ _04291_ VGND VGND VPWR
+ VPWR _00540_ sky130_fd_sc_hd__o211a_1
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11087_ _04784_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__inv_2
Xinput250 hash[94] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_4
X_10038_ sha256cu.msg_scheduler.mreg_1\[19\] _04247_ _04257_ _04250_ VGND VGND VPWR
+ VPWR _00511_ sky130_fd_sc_hd__o211a_1
XFILLER_49_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14915_ clknet_leaf_99_clk _01429_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14846_ clknet_leaf_115_clk _01360_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14777_ clknet_leaf_121_clk _01291_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11989_ _05803_ _05804_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__nor2_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13728_ clknet_leaf_84_clk _00274_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13659_ clknet_leaf_67_clk _00205_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07180_ _00457_ _01843_ _01845_ _01847_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a31o_1
XFILLER_129_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09821_ sha256cu.msg_scheduler.mreg_13\[31\] _04126_ _04131_ _04130_ VGND VGND VPWR
+ VPWR _00414_ sky130_fd_sc_hd__o211a_1
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09752_ sha256cu.msg_scheduler.mreg_14\[2\] _04080_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__or2_1
XFILLER_86_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08703_ _03202_ _03203_ _03204_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__o21ai_1
X_06964_ _01639_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09683_ sha256cu.msg_scheduler.mreg_14\[4\] _04045_ _04052_ _04050_ VGND VGND VPWR
+ VPWR _00355_ sky130_fd_sc_hd__o211a_1
XFILLER_67_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06895_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkinv_2
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08634_ _02923_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__clkbuf_8
XFILLER_66_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08565_ sha256cu.m_out_digest.b_in\[31\] sha256cu.m_out_digest.a_in\[31\] sha256cu.m_out_digest.c_in\[31\]
+ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__a21o_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07516_ _02140_ _02142_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__xor2_2
XFILLER_70_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08496_ _03095_ _03096_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__or2_1
X_07447_ sha256cu.m_out_digest.g_in\[2\] sha256cu.m_out_digest.f_in\[2\] sha256cu.m_out_digest.e_in\[2\]
+ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__mux2_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07378_ sha256cu.counter_iteration\[0\] sha256cu.m_out_digest.temp_delay _02008_
+ _02011_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__or4_1
XFILLER_7_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09117_ _03601_ _03602_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__xor2_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09048_ _02525_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__xor2_1
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11010_ sha256cu.m_pad_pars.block_512\[59\]\[4\] _04829_ _04833_ sha256cu.m_pad_pars.block_512\[55\]\[4\]
+ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a22o_1
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12961_ sha256cu.m_pad_pars.block_512\[35\]\[6\] _06462_ VGND VGND VPWR VPWR _06469_
+ sky130_fd_sc_hd__and2_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ sha256cu.msg_scheduler.mreg_9\[14\] sha256cu.msg_scheduler.mreg_0\[14\] VGND
+ VGND VPWR VPWR _05731_ sky130_fd_sc_hd__or2_1
XANTENNA_300 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14700_ clknet_leaf_7_clk _01214_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12892_ sha256cu.m_pad_pars.block_512\[31\]\[6\] _06425_ VGND VGND VPWR VPWR _06432_
+ sky130_fd_sc_hd__and2_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_311 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11843_ sha256cu.iter_processing.w\[10\] _05430_ _05665_ _05640_ VGND VGND VPWR VPWR
+ _00908_ sky130_fd_sc_hd__o211a_1
XANTENNA_333 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_322 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14631_ clknet_leaf_13_clk _01145_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[26\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_377 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 net207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_366 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_344 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_399 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ sha256cu.msg_scheduler.mreg_9\[8\] sha256cu.msg_scheduler.mreg_0\[8\] VGND
+ VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nand2_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14562_ clknet_leaf_96_clk _01076_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ sha256cu.msg_scheduler.mreg_11\[26\] _04640_ VGND VGND VPWR VPWR _04650_
+ sky130_fd_sc_hd__or2_1
X_14493_ clknet_leaf_121_clk _01007_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13513_ sha256cu.K\[30\] _06716_ _06717_ _06772_ _06737_ VGND VGND VPWR VPWR _01471_
+ sky130_fd_sc_hd__o221a_1
X_10656_ sha256cu.msg_scheduler.mreg_10\[28\] _04601_ VGND VGND VPWR VPWR _04611_
+ sky130_fd_sc_hd__or2_1
X_13444_ sha256cu.K\[4\] _06726_ _06727_ _06729_ _05040_ VGND VGND VPWR VPWR _01445_
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10587_ sha256cu.msg_scheduler.mreg_8\[30\] _04567_ _04571_ _04570_ VGND VGND VPWR
+ VPWR _00746_ sky130_fd_sc_hd__o211a_1
X_13375_ _06688_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_1
X_12326_ _06109_ _06112_ _06126_ _05465_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__a31o_1
XFILLER_141_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12257_ _06059_ _06061_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__xor2_1
XFILLER_141_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12188_ _05994_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__or2_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11208_ sha256cu.m_pad_pars.block_512\[62\]\[5\] _04984_ _04982_ sha256cu.m_pad_pars.block_512\[58\]\[5\]
+ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_150_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11139_ _04768_ _04994_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__nor2_1
XFILLER_64_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14829_ clknet_leaf_8_clk _01343_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08350_ _02953_ _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07301_ sha256cu.byte_stop _01916_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__nand2_2
XFILLER_149_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08281_ sha256cu.K\[23\] _02870_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__and2_1
X_07232_ _01665_ _01648_ _01809_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__and3_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07163_ _01832_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__inv_1
XFILLER_145_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07094_ _01605_ _01647_ _01650_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ sha256cu.msg_scheduler.mreg_14\[24\] _04120_ VGND VGND VPWR VPWR _04122_
+ sky130_fd_sc_hd__or2_1
XFILLER_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07996_ _02563_ _02573_ _02609_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__o21ba_1
XFILLER_86_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09735_ sha256cu.msg_scheduler.mreg_14\[26\] _04073_ _04082_ _04077_ VGND VGND VPWR
+ VPWR _00377_ sky130_fd_sc_hd__o211a_1
XFILLER_55_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06947_ _00452_ _00453_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__or2_2
X_09666_ sha256cu.m_out_digest.h_in\[30\] _02369_ _02478_ sha256cu.m_out_digest.g_in\[30\]
+ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__o22a_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08617_ sha256cu.m_out_digest.c_in\[1\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[1\]
+ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__o22a_1
XFILLER_82_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06878_ sha256cu.counter_iteration\[2\] sha256cu.msg_scheduler.counter_iteration\[2\]
+ _01568_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__mux2_2
X_09597_ _02923_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__buf_4
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08548_ _02304_ _02220_ _03145_ _03147_ _02258_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__a221o_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08479_ sha256cu.m_out_digest.h_in\[29\] _03079_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__xnor2_1
X_10510_ sha256cu.msg_scheduler.mreg_8\[30\] _04520_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__or2_1
X_11490_ sha256cu.m_pad_pars.block_512\[40\]\[1\] _05320_ _05299_ sha256cu.m_pad_pars.block_512\[12\]\[1\]
+ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__a221o_1
XFILLER_11_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10441_ sha256cu.msg_scheduler.mreg_8\[0\] _04481_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__or2_1
XFILLER_109_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10372_ sha256cu.msg_scheduler.mreg_7\[2\] _04441_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__or2_1
X_13160_ sha256cu.m_pad_pars.block_512\[47\]\[3\] _06571_ VGND VGND VPWR VPWR _06575_
+ sky130_fd_sc_hd__and2_1
X_12111_ _05895_ _05899_ _05896_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__a21boi_1
X_13091_ sha256cu.m_pad_pars.block_512\[43\]\[3\] _06534_ VGND VGND VPWR VPWR _06538_
+ sky130_fd_sc_hd__and2_1
X_12042_ sha256cu.msg_scheduler.mreg_14\[29\] _05855_ VGND VGND VPWR VPWR _05856_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13993_ clknet_leaf_57_clk _00539_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12944_ sha256cu.m_pad_pars.block_512\[34\]\[6\] _06453_ VGND VGND VPWR VPWR _06460_
+ sky130_fd_sc_hd__and2_1
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ sha256cu.m_pad_pars.block_512\[30\]\[6\] _06416_ VGND VGND VPWR VPWR _06423_
+ sky130_fd_sc_hd__and2_1
XFILLER_61_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_141 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _05647_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__or2_1
XANTENNA_185 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14614_ clknet_leaf_113_clk _01128_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11757_ _05555_ _05556_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__or2_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14545_ clknet_leaf_7_clk _01059_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_196 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10708_ _04547_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__clkbuf_2
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11688_ _05515_ _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__and2_1
X_14476_ clknet_leaf_8_clk _00990_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10639_ _04547_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__clkbuf_2
X_13427_ sha256cu.iter_processing.padding_done _06716_ VGND VGND VPWR VPWR _06717_
+ sky130_fd_sc_hd__nand2_2
XFILLER_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13358_ _06679_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12309_ _06072_ _06075_ _06090_ _06091_ _06111_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__o311ai_4
XFILLER_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13289_ _06643_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07850_ _02430_ _02432_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__nor2_1
XFILLER_57_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07781_ _02398_ _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__xnor2_1
X_06801_ net235 net238 net237 net240 VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__or4_1
X_09520_ _03990_ _03991_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand2_1
Xinput3 hash[101] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09451_ _03892_ _03921_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__nand2_1
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08402_ _03002_ _03004_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__xor2_1
X_09382_ _03820_ _03824_ _03818_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__o21a_1
X_08333_ sha256cu.m_out_digest.b_in\[25\] sha256cu.m_out_digest.a_in\[25\] _02937_
+ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_125_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_16
X_08264_ sha256cu.K\[23\] _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__xnor2_2
XFILLER_119_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08195_ sha256cu.m_out_digest.a_in\[21\] _02440_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__or2_1
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07215_ _01618_ _01877_ _01679_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07146_ _01710_ _01687_ _01714_ _01621_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__a211o_1
XFILLER_105_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07077_ _01632_ _01615_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__or2_1
XFILLER_105_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07979_ sha256cu.m_out_digest.b_in\[16\] _02128_ sha256cu.m_out_digest.c_in\[16\]
+ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__a21o_1
X_09718_ sha256cu.msg_scheduler.mreg_14\[19\] _04060_ _04072_ _04064_ VGND VGND VPWR
+ VPWR _00370_ sky130_fd_sc_hd__o211a_1
XFILLER_74_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10990_ sha256cu.m_pad_pars.block_512\[39\]\[2\] _04800_ _04831_ sha256cu.m_pad_pars.block_512\[19\]\[2\]
+ _04854_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__a221o_1
X_09649_ sha256cu.m_out_digest.h_in\[13\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[13\]
+ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__a22o_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12660_ sha256cu.m_pad_pars.block_512\[18\]\[1\] _06307_ VGND VGND VPWR VPWR _06309_
+ sky130_fd_sc_hd__and2_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11611_ _05439_ _05441_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__nand2_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _06272_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__clkbuf_1
X_14330_ clknet_leaf_10_clk _00844_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.m_size\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11542_ sha256cu.m_pad_pars.block_512\[44\]\[6\] _05298_ _05304_ sha256cu.m_pad_pars.block_512\[36\]\[6\]
+ _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__a221o_1
XFILLER_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14261_ clknet_leaf_27_clk _00807_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11473_ sha256cu.m_pad_pars.add_512_block\[6\] _04770_ VGND VGND VPWR VPWR _05316_
+ sky130_fd_sc_hd__nor2_1
X_10424_ sha256cu.msg_scheduler.mreg_6\[24\] _04474_ _04478_ _04477_ VGND VGND VPWR
+ VPWR _00676_ sky130_fd_sc_hd__o211a_1
X_14192_ clknet_leaf_29_clk _00738_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_13212_ sha256cu.m_pad_pars.block_512\[50\]\[3\] _06599_ VGND VGND VPWR VPWR _06603_
+ sky130_fd_sc_hd__and2_1
XFILLER_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13143_ sha256cu.m_pad_pars.block_512\[46\]\[3\] _06562_ VGND VGND VPWR VPWR _06566_
+ sky130_fd_sc_hd__and2_1
XFILLER_140_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10355_ sha256cu.msg_scheduler.mreg_6\[27\] _04428_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__or2_1
XFILLER_124_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ sha256cu.msg_scheduler.mreg_4\[29\] _04393_ _04399_ _04397_ VGND VGND VPWR
+ VPWR _00617_ sky130_fd_sc_hd__o211a_1
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13074_ sha256cu.m_pad_pars.block_512\[42\]\[3\] _06525_ VGND VGND VPWR VPWR _06529_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12025_ _05838_ _05839_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__nand2_1
XFILLER_66_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13976_ clknet_leaf_42_clk _00522_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[30\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_46_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12927_ sha256cu.m_pad_pars.block_512\[33\]\[6\] _06444_ VGND VGND VPWR VPWR _06451_
+ sky130_fd_sc_hd__and2_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12858_ sha256cu.m_pad_pars.block_512\[29\]\[6\] _06407_ VGND VGND VPWR VPWR _06414_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _05630_ _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__xnor2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_16
X_12789_ _06377_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14528_ clknet_leaf_106_clk _01042_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14459_ clknet_leaf_126_clk _00973_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07000_ _01604_ _01684_ _01685_ _01585_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__a211o_1
XFILLER_127_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08951_ _03441_ _03442_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__and2_1
XFILLER_130_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08882_ _03374_ _03375_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__or2_1
X_07902_ sha256cu.iter_processing.w\[13\] _02489_ _02517_ VGND VGND VPWR VPWR _02518_
+ sky130_fd_sc_hd__a21o_1
XFILLER_97_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07833_ _02450_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__inv_2
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07764_ sha256cu.m_out_digest.a_in\[23\] _02383_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__xnor2_2
XFILLER_84_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07695_ _02283_ _02281_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__or2b_1
XFILLER_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09503_ sha256cu.K\[28\] _03939_ _03938_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__a21o_1
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09434_ sha256cu.iter_processing.w\[27\] _03008_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__and2_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09365_ _03828_ _03829_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nand2_1
XFILLER_21_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_30 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _03774_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__xnor2_1
X_08316_ _02885_ _02920_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__nand2_1
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_74 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08247_ sha256cu.m_out_digest.h_in\[22\] _02808_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__and2_1
XANTENNA_63 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_85 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08178_ sha256cu.iter_processing.w\[21\] _02786_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__xor2_1
X_07129_ _01631_ _01800_ _01801_ _01803_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__o22a_1
X_10140_ sha256cu.msg_scheduler.mreg_2\[30\] _04315_ _04316_ _04304_ VGND VGND VPWR
+ VPWR _00554_ sky130_fd_sc_hd__o211a_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10071_ _04263_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__buf_2
XFILLER_88_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13830_ clknet_leaf_76_clk _00376_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[25\]
+ sky130_fd_sc_hd__dfxtp_2
X_13761_ clknet_leaf_84_clk _00307_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10973_ sha256cu.data_in_padd\[0\] _04741_ _04742_ _04839_ VGND VGND VPWR VPWR _00863_
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12712_ _06336_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__clkbuf_1
X_13692_ clknet_leaf_67_clk _00238_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[15\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12643_ sha256cu.m_pad_pars.block_512\[17\]\[1\] _06298_ VGND VGND VPWR VPWR _06300_
+ sky130_fd_sc_hd__and2_1
XFILLER_30_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12574_ sha256cu.m_pad_pars.block_512\[13\]\[1\] _06261_ VGND VGND VPWR VPWR _06263_
+ sky130_fd_sc_hd__and2_1
XFILLER_129_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11525_ sha256cu.m_pad_pars.block_512\[0\]\[4\] _05314_ _05360_ _05363_ VGND VGND
+ VPWR VPWR _05364_ sky130_fd_sc_hd__a211o_1
X_14313_ clknet_leaf_91_clk _00006_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__dfxtp_1
X_14244_ clknet_leaf_28_clk _00790_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11456_ _04769_ _05295_ _01936_ _01992_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__o211a_2
X_10407_ sha256cu.msg_scheduler.mreg_7\[17\] _04468_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__or2_1
XFILLER_125_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14175_ clknet_leaf_35_clk _00721_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11387_ _04794_ _04960_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__nor2_1
XFILLER_152_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10338_ sha256cu.msg_scheduler.mreg_5\[19\] _04421_ _04429_ _04424_ VGND VGND VPWR
+ VPWR _00639_ sky130_fd_sc_hd__o211a_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13126_ sha256cu.m_pad_pars.block_512\[45\]\[3\] _06553_ VGND VGND VPWR VPWR _06557_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ sha256cu.m_pad_pars.block_512\[41\]\[3\] _06516_ VGND VGND VPWR VPWR _06520_
+ sky130_fd_sc_hd__and2_1
X_10269_ sha256cu.msg_scheduler.mreg_4\[22\] _04380_ _04389_ _04383_ VGND VGND VPWR
+ VPWR _00610_ sky130_fd_sc_hd__o211a_1
X_12008_ _05821_ _05822_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__nand2_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13959_ clknet_leaf_58_clk _00505_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_94_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07480_ _01564_ _02064_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__nand2_2
XFILLER_148_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09150_ _03615_ _03616_ _03634_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__and3_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09081_ _03566_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__or2_1
X_08101_ sha256cu.m_out_digest.e_in\[30\] _02711_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__xnor2_2
X_08032_ _02233_ sha256cu.m_out_digest.a_in\[7\] VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__xnor2_1
Xinput50 hash[144] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
Xinput61 hash[154] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput72 hash[164] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
Xinput94 hash[184] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
XFILLER_143_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput83 hash[174] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
XFILLER_143_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09983_ sha256cu.msg_scheduler.mreg_0\[27\] _04221_ _04226_ _04224_ VGND VGND VPWR
+ VPWR _00487_ sky130_fd_sc_hd__o211a_1
XFILLER_107_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08934_ _02380_ _03425_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__xor2_1
XFILLER_131_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08865_ _03329_ _03341_ _03359_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__and3_1
XFILLER_85_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07816_ _02409_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__xor2_2
X_08796_ _03291_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__nor2_1
XFILLER_85_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07747_ _02069_ _02367_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__nor2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07678_ sha256cu.iter_processing.w\[8\] _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__xnor2_2
XFILLER_53_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09417_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__inv_2
XFILLER_139_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09348_ _03791_ _03799_ _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__o21ai_1
X_09279_ _03757_ _03758_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__nand2_1
XFILLER_21_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11310_ _01950_ _04704_ _05159_ _05149_ _05152_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__o311a_2
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12290_ _06072_ _06075_ _06092_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__or3_1
X_11241_ sha256cu.m_pad_pars.block_512\[10\]\[7\] _05090_ _05091_ _05092_ VGND VGND
+ VPWR VPWR _05093_ sky130_fd_sc_hd__o211a_1
X_11172_ sha256cu.data_in_padd\[9\] _04741_ _04742_ _05029_ VGND VGND VPWR VPWR _00872_
+ sky130_fd_sc_hd__a22o_1
X_10123_ sha256cu.msg_scheduler.mreg_2\[23\] _04301_ _04306_ _04304_ VGND VGND VPWR
+ VPWR _00547_ sky130_fd_sc_hd__o211a_1
XFILLER_134_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10054_ sha256cu.msg_scheduler.mreg_2\[26\] _04254_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__or2_1
XFILLER_75_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14931_ clknet_leaf_89_clk _01445_ VGND VGND VPWR VPWR sha256cu.K\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14862_ clknet_leaf_11_clk _01376_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13813_ clknet_leaf_49_clk _00359_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14793_ clknet_leaf_13_clk _01307_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13744_ clknet_leaf_66_clk _00290_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10956_ _01952_ _04759_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__nor2_2
X_13675_ clknet_leaf_71_clk _00221_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10887_ _04702_ _04751_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__o21a_1
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12626_ sha256cu.m_pad_pars.block_512\[16\]\[1\] _06289_ VGND VGND VPWR VPWR _06291_
+ sky130_fd_sc_hd__and2_1
XFILLER_129_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12557_ sha256cu.m_pad_pars.block_512\[12\]\[1\] _06252_ VGND VGND VPWR VPWR _06254_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12488_ _06216_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
X_11508_ sha256cu.m_pad_pars.block_512\[4\]\[3\] _05313_ _05320_ sha256cu.m_pad_pars.block_512\[40\]\[3\]
+ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__a22o_1
X_14227_ clknet_leaf_26_clk _00773_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11439_ _04807_ _05136_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__nor2_1
X_14158_ clknet_leaf_31_clk _00704_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ sha256cu.m_pad_pars.block_512\[44\]\[3\] _06544_ VGND VGND VPWR VPWR _06548_
+ sky130_fd_sc_hd__and2_1
X_14089_ clknet_leaf_37_clk _00635_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _01667_ _01634_ _01591_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__o21a_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ sha256cu.m_out_digest.c_in\[30\] _03184_ _03182_ sha256cu.m_out_digest.b_in\[30\]
+ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__a22o_1
X_07601_ _02222_ _02223_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__and3_1
XFILLER_82_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08581_ sha256cu.m_out_digest.b_in\[3\] _03031_ _02114_ sha256cu.m_out_digest.a_in\[3\]
+ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__a22o_1
XFILLER_82_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07532_ sha256cu.m_out_digest.e_in\[15\] sha256cu.m_out_digest.e_in\[10\] VGND VGND
+ VPWR VPWR _02158_ sky130_fd_sc_hd__xnor2_1
X_07463_ _02088_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09202_ _03670_ _03654_ _03683_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__nor3_1
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07394_ sha256cu.m_out_digest.e_in\[25\] _02023_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__xnor2_2
X_09133_ sha256cu.m_out_digest.h_in\[17\] sha256cu.m_out_digest.d_in\[17\] VGND VGND
+ VPWR VPWR _03618_ sky130_fd_sc_hd__nand2_1
XFILLER_135_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09064_ _03520_ _03531_ _03550_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__nand3_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08015_ _02037_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__buf_4
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09966_ sha256cu.msg_scheduler.mreg_1\[20\] _04215_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__or2_1
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08917_ _03408_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__xnor2_1
X_09897_ sha256cu.msg_scheduler.mreg_12\[31\] _04167_ _04175_ _04171_ VGND VGND VPWR
+ VPWR _00446_ sky130_fd_sc_hd__o211a_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _03325_ _03326_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__nor2_1
XFILLER_85_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08779_ _03248_ _03249_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__or2_1
XFILLER_72_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10810_ sha256cu.msg_scheduler.mreg_11\[31\] _04685_ _04697_ _04688_ VGND VGND VPWR
+ VPWR _00843_ sky130_fd_sc_hd__o211a_1
X_11790_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__inv_2
XFILLER_72_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10741_ sha256cu.msg_scheduler.mreg_11\[1\] _04646_ _04658_ _04649_ VGND VGND VPWR
+ VPWR _00813_ sky130_fd_sc_hd__o211a_1
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13460_ sha256cu.K\[10\] _06726_ _06727_ _06739_ _06737_ VGND VGND VPWR VPWR _01451_
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10672_ sha256cu.msg_scheduler.mreg_10\[3\] _04607_ _04619_ _04610_ VGND VGND VPWR
+ VPWR _00783_ sky130_fd_sc_hd__o211a_1
X_12411_ _06175_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
X_13391_ sha256cu.m_pad_pars.block_512\[61\]\[0\] _06693_ VGND VGND VPWR VPWR _06697_
+ sky130_fd_sc_hd__and2_1
X_12342_ sha256cu.m_pad_pars.add_512_block\[4\] _06136_ VGND VGND VPWR VPWR _06139_
+ sky130_fd_sc_hd__or2_1
XFILLER_5_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12273_ _05448_ _06075_ _06076_ _06077_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__o31ai_1
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14012_ clknet_leaf_41_clk _00558_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11224_ sha256cu.m_pad_pars.block_512\[50\]\[6\] _05008_ _05072_ _05076_ VGND VGND
+ VPWR VPWR _05077_ sky130_fd_sc_hd__a211o_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11155_ _04747_ _04994_ _04990_ _04726_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__o211a_2
X_10106_ sha256cu.msg_scheduler.mreg_3\[16\] _04295_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__or2_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11086_ _04753_ _04933_ _04788_ sha256cu.m_pad_pars.block_512\[11\]\[7\] VGND VGND
+ VPWR VPWR _04946_ sky130_fd_sc_hd__o22a_1
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput240 hash[85] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_2
X_10037_ sha256cu.msg_scheduler.mreg_2\[19\] _04254_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__or2_1
Xinput251 hash[95] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_2
XFILLER_64_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_87_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_49_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14914_ clknet_leaf_101_clk _01428_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14845_ clknet_leaf_119_clk _01359_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11988_ _05776_ _05780_ _05777_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__a21boi_1
XFILLER_91_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14776_ clknet_leaf_122_clk _01290_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13727_ clknet_leaf_69_clk _00273_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10939_ sha256cu.m_pad_pars.temp_chk _04744_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__or2_1
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13658_ clknet_leaf_67_clk _00204_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13589_ clknet_leaf_61_clk _00135_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_11_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
X_12609_ sha256cu.m_pad_pars.block_512\[15\]\[1\] _06280_ VGND VGND VPWR VPWR _06282_
+ sky130_fd_sc_hd__and2_1
XFILLER_144_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09820_ sha256cu.msg_scheduler.mreg_14\[31\] _04120_ VGND VGND VPWR VPWR _04131_
+ sky130_fd_sc_hd__or2_1
XFILLER_113_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09751_ sha256cu.msg_scheduler.mreg_13\[1\] _04086_ _04091_ _04090_ VGND VGND VPWR
+ VPWR _00384_ sky130_fd_sc_hd__o211a_1
X_06963_ _01652_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08702_ sha256cu.m_out_digest.e_in\[0\] _02732_ _01913_ VGND VGND VPWR VPWR _03204_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_79_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_78_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09682_ sha256cu.iter_processing.w\[4\] _04046_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__or2_1
XFILLER_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06894_ _01564_ _01587_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__nand2_4
X_08633_ sha256cu.m_out_digest.c_in\[15\] _03181_ _03183_ sha256cu.m_out_digest.b_in\[15\]
+ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__o22a_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08564_ _02382_ sha256cu.m_out_digest.a_in\[1\] VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__xor2_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07515_ _02072_ _02095_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__a21oi_2
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08495_ _03077_ _03055_ _03094_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__and3_1
X_07446_ sha256cu.m_out_digest.b_in\[2\] sha256cu.m_out_digest.a_in\[2\] sha256cu.m_out_digest.c_in\[2\]
+ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__a21o_1
X_07377_ sha256cu.m_out_digest.h_in\[0\] sha256cu.m_out_digest.H7\[0\] VGND VGND VPWR
+ VPWR _02011_ sky130_fd_sc_hd__xor2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09116_ sha256cu.K\[15\] _03569_ _03570_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__a21o_1
X_09047_ _03533_ _03534_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__nand2_1
XFILLER_132_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09949_ sha256cu.msg_scheduler.mreg_1\[13\] _04202_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__or2_1
XFILLER_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12960_ _06468_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ sha256cu.iter_processing.w\[13\] _05666_ _05730_ _05640_ VGND VGND VPWR VPWR
+ _00911_ sky130_fd_sc_hd__o211a_1
XANTENNA_301 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12891_ _06431_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_323 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_334 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ sha256cu.data_in_padd\[10\] _05433_ _05662_ _05664_ _04046_ VGND VGND VPWR
+ VPWR _05665_ sky130_fd_sc_hd__a221o_1
XFILLER_72_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14630_ clknet_leaf_116_clk _01144_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_345 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_356 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_367 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14561_ clknet_leaf_96_clk _01075_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ sha256cu.msg_scheduler.mreg_9\[8\] sha256cu.msg_scheduler.mreg_0\[8\] VGND
+ VGND VPWR VPWR _05598_ sky130_fd_sc_hd__or2_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_378 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_389 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13512_ sha256cu.counter_iteration\[6\] _00059_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__and2b_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ sha256cu.msg_scheduler.mreg_10\[25\] _04646_ _04648_ _04649_ VGND VGND VPWR
+ VPWR _00805_ sky130_fd_sc_hd__o211a_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14492_ clknet_leaf_122_clk _01006_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10655_ sha256cu.msg_scheduler.mreg_9\[27\] _04607_ _04609_ _04610_ VGND VGND VPWR
+ VPWR _00775_ sky130_fd_sc_hd__o211a_1
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13443_ _04188_ _00062_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__and2b_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13374_ sha256cu.m_pad_pars.block_512\[60\]\[0\] _06682_ VGND VGND VPWR VPWR _06688_
+ sky130_fd_sc_hd__and2_1
XFILLER_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10586_ sha256cu.msg_scheduler.mreg_9\[30\] _04561_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__or2_1
X_12325_ _06109_ _06112_ _06126_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12256_ sha256cu.msg_scheduler.mreg_1\[31\] _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12187_ _05968_ _05972_ _05969_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__a21boi_1
X_11207_ sha256cu.m_pad_pars.block_512\[26\]\[5\] _04964_ _05014_ sha256cu.m_pad_pars.block_512\[18\]\[5\]
+ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__a22o_1
XFILLER_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11138_ _04725_ _04721_ sha256cu.m_pad_pars.add_out2\[3\] sha256cu.m_pad_pars.add_out2\[2\]
+ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__or4_2
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
X_11069_ _04766_ _04767_ _04923_ _04928_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__a31o_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14828_ clknet_leaf_7_clk _01342_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14759_ clknet_leaf_8_clk _01273_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07300_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__clkinv_2
X_08280_ _02868_ _02869_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__and2b_1
X_07231_ _01621_ _01615_ _01890_ _01663_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__a31o_1
X_07162_ _01583_ _01830_ _01674_ _01738_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__o32a_1
XFILLER_20_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07093_ _01690_ _01625_ _01603_ _01682_ _01654_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__a32o_1
XFILLER_132_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09803_ sha256cu.msg_scheduler.mreg_13\[23\] _04112_ _04121_ _04117_ VGND VGND VPWR
+ VPWR _00406_ sky130_fd_sc_hd__o211a_1
X_07995_ _02570_ _02572_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nor2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09734_ sha256cu.iter_processing.w\[26\] _04080_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__or2_1
X_06946_ _01590_ _01634_ _01635_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__and3_1
X_09665_ sha256cu.m_out_digest.h_in\[29\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[29\]
+ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__a22o_1
X_06877_ _01571_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_4
X_08616_ _02369_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__buf_4
XFILLER_55_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09596_ sha256cu.m_out_digest.g_in\[1\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[1\]
+ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__o22a_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08547_ _03144_ _03146_ _02069_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__a21oi_1
X_08478_ sha256cu.m_out_digest.a_in\[31\] _03078_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__xnor2_2
X_07429_ _02025_ _02030_ _02057_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__o21a_1
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10440_ _04447_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__buf_2
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10371_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__buf_2
X_12110_ _05918_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__xor2_1
X_13090_ _06537_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12041_ sha256cu.msg_scheduler.mreg_14\[6\] sha256cu.msg_scheduler.mreg_14\[4\] VGND
+ VGND VPWR VPWR _05855_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13992_ clknet_leaf_58_clk _00538_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12943_ _06459_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12874_ _06422_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_142 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_120 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_164 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11825_ _05621_ _05625_ _05622_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__a21boi_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14613_ clknet_leaf_0_clk _01127_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11756_ _05579_ _05581_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__xnor2_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ clknet_leaf_6_clk _01058_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_197 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10707_ sha256cu.msg_scheduler.mreg_10\[18\] _04633_ _04639_ _04636_ VGND VGND VPWR
+ VPWR _00798_ sky130_fd_sc_hd__o211a_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ clknet_leaf_9_clk _00989_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11687_ _05513_ _05514_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__nand2_1
X_13426_ _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__clkbuf_2
X_10638_ sha256cu.msg_scheduler.mreg_9\[20\] _04594_ _04600_ _04597_ VGND VGND VPWR
+ VPWR _00768_ sky130_fd_sc_hd__o211a_1
XFILLER_10_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10569_ _04547_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__clkbuf_2
X_13357_ sha256cu.m_pad_pars.block_512\[59\]\[0\] _06671_ VGND VGND VPWR VPWR _06679_
+ sky130_fd_sc_hd__and2_1
XFILLER_115_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12308_ _06109_ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__and2_1
X_13288_ sha256cu.m_pad_pars.block_512\[54\]\[7\] _05104_ _01965_ VGND VGND VPWR VPWR
+ _06643_ sky130_fd_sc_hd__mux2_1
XFILLER_6_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12239_ _06017_ _06021_ _06044_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__nand3_1
XFILLER_130_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07780_ sha256cu.K\[9\] _02360_ _02399_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__a21oi_1
X_06800_ net226 net229 net228 net231 VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__or4_2
Xinput4 hash[102] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09450_ _02220_ _03922_ _03923_ _03924_ _01984_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__o311a_1
X_08401_ sha256cu.m_out_digest.h_in\[26\] _02961_ _03003_ VGND VGND VPWR VPWR _03004_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_52_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09381_ _03856_ _03857_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__nor2_1
X_08332_ sha256cu.m_out_digest.b_in\[25\] sha256cu.m_out_digest.a_in\[25\] sha256cu.m_out_digest.c_in\[25\]
+ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__a21o_1
XFILLER_20_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08263_ _02868_ _02869_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07214_ _01690_ _01687_ _01609_ _01685_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__a31o_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08194_ _02801_ _02802_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__xor2_1
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07145_ _00455_ _01739_ _01798_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__a21o_1
X_07076_ _01648_ _01687_ _01628_ _01585_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__a211o_1
XFILLER_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07978_ sha256cu.iter_processing.w\[15\] _02562_ _02591_ VGND VGND VPWR VPWR _02592_
+ sky130_fd_sc_hd__a21o_1
XFILLER_101_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09717_ sha256cu.iter_processing.w\[19\] _04067_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__or2_1
XFILLER_68_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06929_ _01596_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__clkbuf_4
X_09648_ sha256cu.m_out_digest.h_in\[12\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[12\]
+ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__a22o_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09579_ sha256cu.m_out_digest.f_in\[19\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[19\]
+ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__a22o_1
XFILLER_55_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11610_ _05439_ _05441_ _05442_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__o21a_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12590_ sha256cu.m_pad_pars.block_512\[14\]\[0\] _06271_ VGND VGND VPWR VPWR _06272_
+ sky130_fd_sc_hd__and2_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11541_ sha256cu.m_pad_pars.block_512\[24\]\[6\] _05279_ _05313_ sha256cu.m_pad_pars.block_512\[4\]\[6\]
+ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__a22o_1
XFILLER_11_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14260_ clknet_leaf_26_clk _00806_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11472_ _01936_ _05278_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__nand2_1
XFILLER_137_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10423_ sha256cu.msg_scheduler.mreg_7\[24\] _04468_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__or2_1
X_14191_ clknet_leaf_31_clk _00737_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13211_ _06602_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_1
X_10354_ sha256cu.msg_scheduler.mreg_5\[26\] _04434_ _04438_ _04437_ VGND VGND VPWR
+ VPWR _00646_ sky130_fd_sc_hd__o211a_1
XFILLER_124_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13142_ _06565_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10285_ sha256cu.msg_scheduler.mreg_5\[29\] _04387_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__or2_1
X_13073_ _06528_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ _05835_ _05836_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__nand2_1
XFILLER_39_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13975_ clknet_leaf_42_clk _00521_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[29\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_65_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12926_ _06450_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__clkbuf_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12857_ _06413_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ sha256cu.msg_scheduler.mreg_14\[28\] _05631_ VGND VGND VPWR VPWR _05632_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_61_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ sha256cu.m_pad_pars.block_512\[25\]\[5\] _06371_ VGND VGND VPWR VPWR _06377_
+ sky130_fd_sc_hd__and2_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11739_ _05525_ _05545_ _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__o21ai_1
X_14527_ clknet_leaf_79_clk _01041_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14458_ clknet_leaf_126_clk _00972_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14389_ clknet_leaf_15_clk _00903_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_13409_ sha256cu.m_pad_pars.m_size\[9\] sha256cu.m_pad_pars.block_512\[62\]\[1\]
+ _01923_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__mux2_1
X_08950_ _03421_ _03422_ _03440_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__nand3_1
X_08881_ _03373_ _03372_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__and2b_1
X_07901_ _02487_ _02488_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__and2b_1
X_07832_ sha256cu.m_out_digest.e_in\[23\] _02449_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__xnor2_2
XFILLER_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07763_ _02382_ sha256cu.m_out_digest.a_in\[0\] VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09502_ _03973_ _03974_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__nor2_1
X_07694_ _02293_ _02315_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__xnor2_2
X_09433_ _03907_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__inv_2
X_09364_ sha256cu.m_out_digest.e_in\[24\] _02732_ _03840_ _03841_ _01913_ VGND VGND
+ VPWR VPWR _00247_ sky130_fd_sc_hd__a221o_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08315_ _02885_ _02920_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__or2_1
XANTENNA_20 _01994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ sha256cu.K\[21\] _03739_ _03738_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__a21o_1
XFILLER_21_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_75 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08246_ sha256cu.m_out_digest.h_in\[22\] _02808_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__or2_1
XANTENNA_64 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_86 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08177_ _02784_ _02785_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__xnor2_1
XANTENNA_97 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07128_ _01631_ _01802_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__nand2_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07059_ _01585_ _01737_ _01738_ _01740_ _01663_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__o311a_1
X_10070_ sha256cu.msg_scheduler.mreg_3\[1\] _04268_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__or2_1
XFILLER_99_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13760_ clknet_leaf_84_clk _00306_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10972_ _04783_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__or2_1
XFILLER_44_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13691_ clknet_leaf_67_clk _00237_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[14\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12711_ sha256cu.m_pad_pars.block_512\[21\]\[1\] _06334_ VGND VGND VPWR VPWR _06336_
+ sky130_fd_sc_hd__and2_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12642_ _06299_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12573_ _06262_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11524_ sha256cu.m_pad_pars.block_512\[52\]\[4\] _05310_ _05288_ sha256cu.m_pad_pars.block_512\[48\]\[4\]
+ _05362_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__a221o_1
XFILLER_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14312_ clknet_leaf_92_clk _00005_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__dfxtp_1
X_14243_ clknet_leaf_28_clk _00789_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11455_ _04912_ _05295_ _05297_ _01992_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__o211a_2
X_10406_ _04414_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__clkbuf_2
XFILLER_109_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14174_ clknet_leaf_45_clk _00720_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11386_ sha256cu.data_in_padd\[22\] _04741_ _04742_ _05230_ VGND VGND VPWR VPWR _00885_
+ sky130_fd_sc_hd__a22o_1
X_10337_ sha256cu.msg_scheduler.mreg_6\[19\] _04428_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__or2_1
X_13125_ _06556_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ sha256cu.msg_scheduler.mreg_5\[22\] _04387_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__or2_1
XFILLER_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13056_ _06519_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__clkbuf_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12007_ sha256cu.msg_scheduler.mreg_9\[18\] sha256cu.msg_scheduler.mreg_0\[18\] VGND
+ VGND VPWR VPWR _05822_ sky130_fd_sc_hd__nand2_1
XFILLER_66_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10199_ sha256cu.msg_scheduler.mreg_4\[24\] _04348_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__or2_1
XFILLER_47_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13958_ clknet_leaf_59_clk _00504_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12909_ sha256cu.m_pad_pars.block_512\[32\]\[6\] _06434_ VGND VGND VPWR VPWR _06441_
+ sky130_fd_sc_hd__and2_1
X_13889_ clknet_leaf_24_clk _00435_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09080_ _03564_ _03565_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__and2_1
X_08100_ sha256cu.m_out_digest.e_in\[25\] sha256cu.m_out_digest.e_in\[12\] VGND VGND
+ VPWR VPWR _02711_ sky130_fd_sc_hd__xnor2_2
X_08031_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__inv_2
Xinput40 hash[135] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
Xinput73 hash[165] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xinput62 hash[155] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
Xinput51 hash[145] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
Xinput95 hash[185] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput84 hash[175] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_143_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09982_ sha256cu.msg_scheduler.mreg_1\[27\] _04215_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__or2_1
X_08933_ _03423_ _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__nand2_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08864_ _03342_ _03358_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07815_ sha256cu.K\[11\] _02433_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__xnor2_2
X_08795_ sha256cu.m_out_digest.h_in\[5\] sha256cu.m_out_digest.d_in\[5\] VGND VGND
+ VPWR VPWR _03292_ sky130_fd_sc_hd__and2_1
XFILLER_96_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07746_ _02364_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07677_ _02297_ _02298_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__and2b_1
X_09416_ _03890_ _03891_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__and2_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09347_ _03820_ _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__xor2_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09278_ sha256cu.m_out_digest.h_in\[22\] sha256cu.m_out_digest.d_in\[22\] VGND VGND
+ VPWR VPWR _03758_ sky130_fd_sc_hd__nand2_1
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08229_ _02805_ _02797_ _02836_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11240_ _04959_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__inv_2
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11171_ sha256cu.m_pad_pars.block_512\[14\]\[1\] _04989_ _05019_ _05028_ VGND VGND
+ VPWR VPWR _05029_ sky130_fd_sc_hd__a211o_1
X_10122_ sha256cu.msg_scheduler.mreg_3\[23\] _04295_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__or2_1
XFILLER_106_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10053_ sha256cu.msg_scheduler.mreg_1\[25\] _04260_ _04266_ _04264_ VGND VGND VPWR
+ VPWR _00517_ sky130_fd_sc_hd__o211a_1
XFILLER_48_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14930_ clknet_leaf_89_clk _01444_ VGND VGND VPWR VPWR sha256cu.K\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14861_ clknet_leaf_11_clk _01375_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13812_ clknet_leaf_47_clk _00358_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_91_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14792_ clknet_leaf_13_clk _01306_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13743_ clknet_leaf_73_clk _00289_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10955_ _04705_ _04820_ _04821_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__o21a_2
X_13674_ clknet_leaf_82_clk _00220_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10886_ _04749_ _04752_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__or2_2
X_12625_ _06290_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12556_ _06253_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__clkbuf_1
X_11507_ sha256cu.m_pad_pars.block_512\[32\]\[3\] _05306_ _05318_ sha256cu.m_pad_pars.block_512\[8\]\[3\]
+ _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__a221o_1
XFILLER_12_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12487_ sha256cu.m_pad_pars.block_512\[8\]\[1\] _06214_ VGND VGND VPWR VPWR _06216_
+ sky130_fd_sc_hd__and2_1
X_14226_ clknet_leaf_26_clk _00772_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[24\]
+ sky130_fd_sc_hd__dfxtp_2
X_11438_ sha256cu.m_pad_pars.block_512\[60\]\[0\] _01998_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[0\]
+ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__a22o_1
X_14157_ clknet_leaf_32_clk _00703_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11369_ sha256cu.m_pad_pars.block_512\[61\]\[5\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[5\]
+ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__a22o_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13108_ _06547_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__clkbuf_1
X_14088_ clknet_leaf_37_clk _00634_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _06510_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07600_ sha256cu.m_out_digest.g_in\[6\] sha256cu.m_out_digest.f_in\[6\] sha256cu.m_out_digest.e_in\[6\]
+ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__mux2_1
X_08580_ sha256cu.m_out_digest.b_in\[2\] _02370_ _02110_ sha256cu.m_out_digest.a_in\[2\]
+ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__o22a_1
XFILLER_82_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07531_ sha256cu.iter_processing.w\[4\] _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07462_ _02052_ _02055_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__o21a_1
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07393_ sha256cu.m_out_digest.e_in\[11\] sha256cu.m_out_digest.e_in\[6\] VGND VGND
+ VPWR VPWR _02023_ sky130_fd_sc_hd__xnor2_1
X_09201_ _03670_ _03654_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__o21a_1
XFILLER_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09132_ sha256cu.m_out_digest.h_in\[17\] sha256cu.m_out_digest.d_in\[17\] VGND VGND
+ VPWR VPWR _03617_ sky130_fd_sc_hd__or2_1
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09063_ _03520_ _03531_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__a21o_1
XFILLER_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08014_ _02621_ _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__nand2_1
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09965_ sha256cu.msg_scheduler.mreg_0\[19\] _04208_ _04216_ _04211_ VGND VGND VPWR
+ VPWR _00479_ sky130_fd_sc_hd__o211a_1
XFILLER_89_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08916_ _03375_ _03381_ _03374_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__o21ba_1
X_09896_ sha256cu.msg_scheduler.mreg_13\[31\] _04174_ VGND VGND VPWR VPWR _04175_
+ sky130_fd_sc_hd__or2_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ sha256cu.K\[6\] _03320_ _03319_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__a21o_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08778_ _03270_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__xor2_1
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07729_ sha256cu.m_out_digest.h_in\[8\] _02306_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__nand2_1
XFILLER_26_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10740_ sha256cu.msg_scheduler.mreg_12\[1\] _04653_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__or2_1
XFILLER_53_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10671_ sha256cu.msg_scheduler.mreg_11\[3\] _04614_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__or2_1
XFILLER_80_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12410_ sha256cu.m_pad_pars.block_512\[3\]\[5\] _06169_ VGND VGND VPWR VPWR _06175_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _06696_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12341_ _06138_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12272_ sha256cu.data_in_padd\[28\] _05433_ _04046_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14011_ clknet_leaf_42_clk _00557_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11223_ sha256cu.m_pad_pars.block_512\[26\]\[6\] _04964_ _05009_ sha256cu.m_pad_pars.block_512\[30\]\[6\]
+ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__a221o_1
XFILLER_5_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11154_ _05011_ _05012_ _04726_ _04951_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__and4bb_2
XFILLER_1_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10105_ sha256cu.msg_scheduler.mreg_2\[15\] _04288_ _04296_ _04291_ VGND VGND VPWR
+ VPWR _00539_ sky130_fd_sc_hd__o211a_1
XFILLER_103_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11085_ sha256cu.m_pad_pars.block_512\[27\]\[7\] _04944_ _04753_ _04907_ VGND VGND
+ VPWR VPWR _04945_ sky130_fd_sc_hd__o22a_1
Xinput230 hash[76] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_2
X_10036_ sha256cu.msg_scheduler.mreg_1\[18\] _04247_ _04256_ _04250_ VGND VGND VPWR
+ VPWR _00510_ sky130_fd_sc_hd__o211a_1
Xinput252 hash[96] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_2
Xinput241 hash[86] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14913_ clknet_leaf_99_clk _01427_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14844_ clknet_leaf_115_clk _01358_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11987_ _05800_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__xor2_1
XFILLER_91_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14775_ clknet_leaf_125_clk _01289_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13726_ clknet_leaf_70_clk _00272_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10938_ sha256cu.m_pad_pars.add_512_block\[6\] _04744_ VGND VGND VPWR VPWR _04805_
+ sky130_fd_sc_hd__or2_1
XFILLER_90_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13657_ clknet_leaf_64_clk _00203_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10869_ _04735_ _04733_ _04739_ _01913_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__a211oi_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13588_ clknet_leaf_59_clk _00134_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12608_ _06281_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__clkbuf_1
X_12539_ _06243_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14209_ clknet_leaf_28_clk _00755_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09750_ sha256cu.msg_scheduler.mreg_14\[1\] _04080_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__or2_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06962_ _01596_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__clkbuf_4
X_09681_ sha256cu.msg_scheduler.mreg_14\[3\] _04045_ _04051_ _04050_ VGND VGND VPWR
+ VPWR _00354_ sky130_fd_sc_hd__o211a_1
X_08701_ _03197_ _03201_ _02629_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__a21o_1
XFILLER_67_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08632_ _02109_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__buf_4
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06893_ sha256cu.counter_iteration\[3\] sha256cu.msg_scheduler.counter_iteration\[3\]
+ _01568_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_82_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08563_ _03153_ _03161_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07514_ _02094_ _02092_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__and2b_1
X_08494_ _03077_ _03055_ _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07445_ sha256cu.m_out_digest.b_in\[2\] sha256cu.m_out_digest.a_in\[2\] VGND VGND
+ VPWR VPWR _02073_ sky130_fd_sc_hd__or2_1
XFILLER_50_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07376_ sha256cu.m_out_digest.temp_delay _02009_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__and2b_1
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09115_ _03599_ _03600_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09046_ sha256cu.m_out_digest.h_in\[14\] sha256cu.m_out_digest.d_in\[14\] VGND VGND
+ VPWR VPWR _03534_ sky130_fd_sc_hd__nand2_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09948_ sha256cu.msg_scheduler.mreg_0\[12\] _04195_ _04206_ _04198_ VGND VGND VPWR
+ VPWR _00472_ sky130_fd_sc_hd__o211a_1
XFILLER_89_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09879_ sha256cu.msg_scheduler.mreg_12\[24\] _04153_ _04164_ _04157_ VGND VGND VPWR
+ VPWR _00439_ sky130_fd_sc_hd__o211a_1
XFILLER_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11910_ sha256cu.data_in_padd\[13\] _05667_ _05729_ _05463_ VGND VGND VPWR VPWR _05730_
+ sky130_fd_sc_hd__a211o_1
X_12890_ sha256cu.m_pad_pars.block_512\[31\]\[5\] _06425_ VGND VGND VPWR VPWR _06431_
+ sky130_fd_sc_hd__and2_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _05660_ _05663_ _05465_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a21oi_1
XANTENNA_324 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_302 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_346 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_368 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_357 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _05583_ _05560_ _05582_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a31o_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14560_ clknet_leaf_96_clk _01074_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _04529_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__buf_2
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13511_ _06771_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ clknet_leaf_121_clk _01005_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10654_ _04529_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__buf_2
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13442_ sha256cu.K\[3\] _06726_ _06727_ _06728_ _05040_ VGND VGND VPWR VPWR _01444_
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10585_ sha256cu.msg_scheduler.mreg_8\[29\] _04567_ _04569_ _04570_ VGND VGND VPWR
+ VPWR _00745_ sky130_fd_sc_hd__o211a_1
X_13373_ _06687_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__clkbuf_1
X_12324_ _06118_ _06125_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12255_ sha256cu.msg_scheduler.mreg_1\[14\] sha256cu.msg_scheduler.mreg_1\[3\] VGND
+ VGND VPWR VPWR _06060_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12186_ _05991_ _05993_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__xor2_1
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11206_ sha256cu.data_in_padd\[12\] _04840_ _05057_ _05060_ _05040_ VGND VGND VPWR
+ VPWR _00875_ sky130_fd_sc_hd__o221a_1
XFILLER_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11137_ _04991_ _04995_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__nor2_4
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11068_ _04756_ _04767_ _04927_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__and3_1
X_10019_ sha256cu.msg_scheduler.mreg_1\[11\] _04234_ _04246_ _04237_ VGND VGND VPWR
+ VPWR _00503_ sky130_fd_sc_hd__o211a_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14827_ clknet_leaf_7_clk _01341_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14758_ clknet_leaf_102_clk _01272_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13709_ clknet_leaf_70_clk _00255_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14689_ clknet_leaf_103_clk _01203_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_07230_ _00454_ _01637_ _01682_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07161_ _01639_ _01696_ _01596_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__a21o_1
XFILLER_117_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07092_ _00457_ _01764_ _01765_ _01770_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__a31o_1
XFILLER_132_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09802_ sha256cu.msg_scheduler.mreg_14\[23\] _04120_ VGND VGND VPWR VPWR _04121_
+ sky130_fd_sc_hd__or2_1
XFILLER_140_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07994_ _02597_ _02607_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__xor2_1
X_09733_ sha256cu.msg_scheduler.mreg_14\[25\] _04073_ _04081_ _04077_ VGND VGND VPWR
+ VPWR _00376_ sky130_fd_sc_hd__o211a_1
X_06945_ _01586_ _01580_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__nand2_1
XFILLER_28_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09664_ sha256cu.m_out_digest.h_in\[28\] _02369_ _02478_ sha256cu.m_out_digest.g_in\[28\]
+ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__o22a_1
XFILLER_27_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06876_ _01570_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__clkinv_2
XFILLER_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09595_ sha256cu.m_out_digest.g_in\[0\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[0\]
+ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__o22a_1
X_08615_ sha256cu.m_out_digest.c_in\[0\] _03179_ _03178_ sha256cu.m_out_digest.b_in\[0\]
+ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__a22o_1
XFILLER_82_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08546_ _03068_ _03071_ _03105_ _03106_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__a31o_1
XFILLER_23_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08477_ _02233_ sha256cu.m_out_digest.a_in\[10\] VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__xnor2_1
X_07428_ sha256cu.m_out_digest.h_in\[0\] _02029_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__nand2_1
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07359_ _01996_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10370_ _04043_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__clkbuf_4
X_09029_ _03512_ _03516_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__and2_1
XFILLER_108_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ _05852_ _05853_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nor2_1
XFILLER_105_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13991_ clknet_leaf_58_clk _00537_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12942_ sha256cu.m_pad_pars.block_512\[34\]\[5\] _06453_ VGND VGND VPWR VPWR _06459_
+ sky130_fd_sc_hd__and2_1
XFILLER_65_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12873_ sha256cu.m_pad_pars.block_512\[30\]\[5\] _06416_ VGND VGND VPWR VPWR _06422_
+ sky130_fd_sc_hd__and2_1
X_14612_ clknet_leaf_5_clk _01126_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_143 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _05644_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__xor2_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_198 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11755_ sha256cu.msg_scheduler.mreg_14\[26\] _05580_ VGND VGND VPWR VPWR _05581_
+ sky130_fd_sc_hd__xnor2_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_187 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14543_ clknet_leaf_6_clk _01057_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10706_ sha256cu.msg_scheduler.mreg_11\[18\] _04627_ VGND VGND VPWR VPWR _04639_
+ sky130_fd_sc_hd__or2_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14474_ clknet_leaf_12_clk _00988_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11686_ _05513_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__or2_1
X_13425_ sha256cu.temp_case _04177_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__or2_1
X_10637_ sha256cu.msg_scheduler.mreg_10\[20\] _04588_ VGND VGND VPWR VPWR _04600_
+ sky130_fd_sc_hd__or2_1
X_10568_ sha256cu.msg_scheduler.mreg_8\[22\] _04554_ _04560_ _04557_ VGND VGND VPWR
+ VPWR _00738_ sky130_fd_sc_hd__o211a_1
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13356_ _06678_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10499_ sha256cu.msg_scheduler.mreg_8\[25\] _04520_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__or2_1
X_12307_ _06107_ _06108_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__nand2_1
X_13287_ _06642_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12238_ _06042_ _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12169_ sha256cu.msg_scheduler.mreg_14\[11\] sha256cu.msg_scheduler.mreg_14\[9\]
+ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__xor2_1
XFILLER_111_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 hash[103] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08400_ _02962_ _02964_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__or2b_1
XFILLER_18_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09380_ _03850_ _03855_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__and2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08331_ _02932_ _02935_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__xor2_1
XFILLER_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08262_ _02829_ _02831_ _02827_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o21bai_1
XFILLER_20_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07213_ _01581_ _01655_ _01618_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__o21a_1
X_08193_ _02758_ _02760_ _02761_ _02767_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__o22a_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07144_ _01812_ _01813_ _01816_ _00457_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__o22a_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07075_ _00455_ _01750_ _01680_ _01715_ _01621_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__a311o_1
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07977_ _02560_ _02561_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__and2b_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09716_ sha256cu.msg_scheduler.mreg_14\[18\] _04060_ _04071_ _04064_ VGND VGND VPWR
+ VPWR _00369_ sky130_fd_sc_hd__o211a_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06928_ _01604_ _01610_ _01616_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__a211o_1
XFILLER_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06859_ net54 net58 net57 net60 VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__or4_1
XFILLER_83_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09647_ _02923_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__clkbuf_4
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09578_ sha256cu.m_out_digest.f_in\[18\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[18\]
+ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__o22a_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08529_ _03123_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__and2_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11540_ sha256cu.m_pad_pars.block_512\[32\]\[6\] _05306_ _05320_ sha256cu.m_pad_pars.block_512\[40\]\[6\]
+ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__a221o_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ _01942_ _04775_ _01937_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__a21oi_4
XFILLER_152_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10422_ sha256cu.msg_scheduler.mreg_6\[23\] _04474_ _04476_ _04477_ VGND VGND VPWR
+ VPWR _00675_ sky130_fd_sc_hd__o211a_1
X_14190_ clknet_leaf_29_clk _00736_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13210_ sha256cu.m_pad_pars.block_512\[50\]\[2\] _06599_ VGND VGND VPWR VPWR _06602_
+ sky130_fd_sc_hd__and2_1
X_10353_ sha256cu.msg_scheduler.mreg_6\[26\] _04428_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__or2_1
X_13141_ sha256cu.m_pad_pars.block_512\[46\]\[2\] _06562_ VGND VGND VPWR VPWR _06565_
+ sky130_fd_sc_hd__and2_1
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13072_ sha256cu.m_pad_pars.block_512\[42\]\[2\] _06525_ VGND VGND VPWR VPWR _06528_
+ sky130_fd_sc_hd__and2_1
X_10284_ sha256cu.msg_scheduler.mreg_4\[28\] _04393_ _04398_ _04397_ VGND VGND VPWR
+ VPWR _00616_ sky130_fd_sc_hd__o211a_1
XFILLER_105_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12023_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__inv_2
XFILLER_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13974_ clknet_leaf_42_clk _00520_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[28\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_93_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12925_ sha256cu.m_pad_pars.block_512\[33\]\[5\] _06444_ VGND VGND VPWR VPWR _06450_
+ sky130_fd_sc_hd__and2_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12856_ sha256cu.m_pad_pars.block_512\[29\]\[5\] _06407_ VGND VGND VPWR VPWR _06413_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ sha256cu.msg_scheduler.mreg_14\[26\] sha256cu.msg_scheduler.mreg_14\[19\]
+ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__xnor2_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _06376_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14526_ clknet_leaf_114_clk _01040_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11738_ _05521_ _05544_ _05543_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__a21o_1
XFILLER_128_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11669_ _05475_ _05477_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__a21oi_1
X_14457_ clknet_leaf_126_clk _00971_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14388_ clknet_leaf_47_clk _00902_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_13408_ _06705_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__clkbuf_1
X_13339_ _06669_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08880_ _03372_ _03373_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__and2b_1
X_07900_ _02027_ _02220_ _02514_ _02516_ _02258_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__a221o_1
X_07831_ sha256cu.m_out_digest.e_in\[18\] sha256cu.m_out_digest.e_in\[5\] VGND VGND
+ VPWR VPWR _02449_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07762_ sha256cu.m_out_digest.a_in\[12\] VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__clkbuf_4
X_09501_ _03934_ _03941_ _03972_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__nor3_1
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07693_ _02312_ _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__xnor2_2
XFILLER_53_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09432_ sha256cu.iter_processing.w\[27\] _03008_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__or2_1
XFILLER_52_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09363_ _03834_ _03839_ _02629_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__a21oi_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08314_ _02918_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__or2b_2
XFILLER_21_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_21 _01994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _01521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09294_ _03772_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__and2_1
XFILLER_21_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_65 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08245_ _02849_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__xnor2_1
XANTENNA_54 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ sha256cu.m_out_digest.g_in\[21\] sha256cu.m_out_digest.f_in\[21\] sha256cu.m_out_digest.e_in\[21\]
+ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__mux2_2
XANTENNA_98 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07127_ _01642_ _01647_ _01594_ _01726_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__a31o_1
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07058_ _01726_ _01739_ _01706_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__or3b_1
XFILLER_153_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10971_ _04813_ _04837_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__or2_1
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13690_ clknet_leaf_64_clk _00236_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_56_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ _06335_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12641_ sha256cu.m_pad_pars.block_512\[17\]\[0\] _06298_ VGND VGND VPWR VPWR _06299_
+ sky130_fd_sc_hd__and2_1
XFILLER_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12572_ sha256cu.m_pad_pars.block_512\[13\]\[0\] _06261_ VGND VGND VPWR VPWR _06262_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14311_ clknet_leaf_93_clk _00004_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11523_ sha256cu.m_pad_pars.block_512\[28\]\[4\] _05296_ _05361_ _01920_ VGND VGND
+ VPWR VPWR _05362_ sky130_fd_sc_hd__a22o_1
X_14242_ clknet_leaf_28_clk _00788_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11454_ sha256cu.m_pad_pars.add_out0\[4\] sha256cu.m_pad_pars.add_out0\[5\] VGND
+ VGND VPWR VPWR _05297_ sky130_fd_sc_hd__nor2b_2
X_10405_ sha256cu.msg_scheduler.mreg_6\[16\] _04461_ _04467_ _04464_ VGND VGND VPWR
+ VPWR _00668_ sky130_fd_sc_hd__o211a_1
X_14173_ clknet_leaf_45_clk _00719_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11385_ sha256cu.m_pad_pars.block_512\[45\]\[6\] _05126_ _05221_ _05229_ VGND VGND
+ VPWR VPWR _05230_ sky130_fd_sc_hd__a211o_1
X_10336_ _04414_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__clkbuf_2
XFILLER_140_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13124_ sha256cu.m_pad_pars.block_512\[45\]\[2\] _06553_ VGND VGND VPWR VPWR _06556_
+ sky130_fd_sc_hd__and2_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ sha256cu.msg_scheduler.mreg_4\[21\] _04380_ _04388_ _04383_ VGND VGND VPWR
+ VPWR _00609_ sky130_fd_sc_hd__o211a_1
XFILLER_112_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_13055_ sha256cu.m_pad_pars.block_512\[41\]\[2\] _06516_ VGND VGND VPWR VPWR _06519_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ sha256cu.msg_scheduler.mreg_9\[18\] sha256cu.msg_scheduler.mreg_0\[18\] VGND
+ VGND VPWR VPWR _05821_ sky130_fd_sc_hd__or2_1
XFILLER_87_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10198_ sha256cu.msg_scheduler.mreg_3\[23\] _04341_ _04349_ _04344_ VGND VGND VPWR
+ VPWR _00579_ sky130_fd_sc_hd__o211a_1
XFILLER_94_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13957_ clknet_leaf_59_clk _00503_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12908_ _06440_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__clkbuf_1
X_13888_ clknet_leaf_24_clk _00434_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ sha256cu.m_pad_pars.block_512\[28\]\[5\] _06398_ VGND VGND VPWR VPWR _06404_
+ sky130_fd_sc_hd__and2_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14509_ clknet_leaf_22_clk _01023_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08030_ sha256cu.m_out_digest.e_in\[28\] _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__xnor2_4
Xinput30 hash[126] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
Xinput52 hash[146] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
Xinput41 hash[136] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput63 hash[156] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xinput85 hash[176] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput74 hash[166] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xinput96 hash[186] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
X_09981_ sha256cu.msg_scheduler.mreg_0\[26\] _04221_ _04225_ _04224_ VGND VGND VPWR
+ VPWR _00486_ sky130_fd_sc_hd__o211a_1
XFILLER_89_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08932_ sha256cu.m_out_digest.h_in\[10\] sha256cu.m_out_digest.d_in\[10\] VGND VGND
+ VPWR VPWR _03424_ sky130_fd_sc_hd__nand2_1
XFILLER_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08863_ _03356_ _03357_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__and2_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07814_ _02430_ _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__xor2_2
X_08794_ sha256cu.m_out_digest.h_in\[5\] sha256cu.m_out_digest.d_in\[5\] VGND VGND
+ VPWR VPWR _03291_ sky130_fd_sc_hd__nor2_1
XFILLER_123_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07745_ _02323_ _02329_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07676_ _02294_ _02295_ _02296_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__a21o_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09415_ _03887_ _03889_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__or2_1
XFILLER_13_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09346_ sha256cu.K\[24\] _03823_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09277_ sha256cu.m_out_digest.h_in\[22\] sha256cu.m_out_digest.d_in\[22\] VGND VGND
+ VPWR VPWR _03757_ sky130_fd_sc_hd__or2_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08228_ _02806_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08159_ _02761_ _02767_ _02478_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__a21o_1
X_11170_ sha256cu.m_pad_pars.block_512\[42\]\[1\] _05001_ _05021_ _05023_ _05027_
+ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__a2111o_1
X_10121_ sha256cu.msg_scheduler.mreg_2\[22\] _04301_ _04305_ _04304_ VGND VGND VPWR
+ VPWR _00546_ sky130_fd_sc_hd__o211a_1
XFILLER_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10052_ sha256cu.msg_scheduler.mreg_2\[25\] _04254_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__or2_1
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14860_ clknet_leaf_7_clk _01374_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13811_ clknet_leaf_49_clk _00357_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_91_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14791_ clknet_leaf_11_clk _01305_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[46\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13742_ clknet_leaf_71_clk _00288_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10954_ _04730_ _04814_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__nor2_1
XFILLER_32_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13673_ clknet_leaf_82_clk _00219_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10885_ _01939_ sha256cu.m_pad_pars.add_512_block\[1\] VGND VGND VPWR VPWR _04752_
+ sky130_fd_sc_hd__or2b_1
X_12624_ sha256cu.m_pad_pars.block_512\[16\]\[0\] _06289_ VGND VGND VPWR VPWR _06290_
+ sky130_fd_sc_hd__and2_1
X_12555_ sha256cu.m_pad_pars.block_512\[12\]\[0\] _06252_ VGND VGND VPWR VPWR _06253_
+ sky130_fd_sc_hd__and2_1
X_11506_ sha256cu.m_pad_pars.block_512\[24\]\[3\] _05279_ _05298_ sha256cu.m_pad_pars.block_512\[44\]\[3\]
+ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__a22o_1
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12486_ _06215_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__clkbuf_1
X_14225_ clknet_leaf_26_clk _00771_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[23\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11437_ sha256cu.m_pad_pars.add_out0\[5\] sha256cu.m_pad_pars.add_out0\[4\] _05278_
+ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__and3_2
XFILLER_153_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14156_ clknet_leaf_32_clk _00702_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11368_ sha256cu.m_pad_pars.block_512\[1\]\[5\] _05135_ _05138_ sha256cu.m_pad_pars.block_512\[17\]\[5\]
+ _05213_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__a221o_1
X_10319_ sha256cu.msg_scheduler.mreg_5\[11\] _04407_ _04418_ _04410_ VGND VGND VPWR
+ VPWR _00631_ sky130_fd_sc_hd__o211a_1
XFILLER_98_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ sha256cu.m_pad_pars.block_512\[44\]\[2\] _06544_ VGND VGND VPWR VPWR _06547_
+ sky130_fd_sc_hd__and2_1
X_14087_ clknet_leaf_38_clk _00633_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _05134_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__and2_1
XFILLER_121_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ sha256cu.m_pad_pars.block_512\[40\]\[2\] _06507_ VGND VGND VPWR VPWR _06510_
+ sky130_fd_sc_hd__and2_1
XFILLER_94_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07530_ _02154_ _02155_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__and2b_1
XFILLER_82_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07461_ sha256cu.m_out_digest.h_in\[1\] _02054_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__nand2_1
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07392_ sha256cu.iter_processing.w\[0\] _02021_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__xnor2_1
X_09200_ _03681_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__nor2_1
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09131_ _03601_ _03602_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__nand2_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09062_ _03548_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08013_ _02623_ _02626_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__and2_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09964_ sha256cu.msg_scheduler.mreg_1\[19\] _04215_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__or2_1
X_08915_ _03403_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__xor2_1
X_09895_ _04133_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__buf_2
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _03331_ _03332_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__nand2_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _03271_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07728_ _02345_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07659_ _02237_ _02239_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__nor2_1
XFILLER_53_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10670_ sha256cu.msg_scheduler.mreg_10\[2\] _04607_ _04618_ _04610_ VGND VGND VPWR
+ VPWR _00782_ sky130_fd_sc_hd__o211a_1
X_09329_ _03772_ _03785_ _03806_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12340_ _06136_ _01983_ _06137_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__and3b_1
X_12271_ _06074_ _06054_ _06056_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__and3_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14010_ clknet_leaf_42_clk _00556_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11222_ sha256cu.m_pad_pars.block_512\[46\]\[6\] _04977_ _04981_ sha256cu.m_pad_pars.block_512\[54\]\[6\]
+ _05074_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__a221o_1
XFILLER_122_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11153_ _04746_ _04954_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__nor2_2
XFILLER_1_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput220 hash[67] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_1
X_10104_ sha256cu.msg_scheduler.mreg_3\[15\] _04295_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__or2_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11084_ _04751_ _04698_ _04908_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__and3b_1
XFILLER_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput231 hash[77] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_2
X_10035_ sha256cu.msg_scheduler.mreg_2\[18\] _04254_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__or2_1
XFILLER_88_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput242 hash[87] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14912_ clknet_leaf_99_clk _01426_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput253 hash[97] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14843_ clknet_leaf_118_clk _01357_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11986_ sha256cu.msg_scheduler.mreg_1\[24\] _05801_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__xnor2_1
X_14774_ clknet_leaf_114_clk _01288_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13725_ clknet_leaf_68_clk _00271_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10937_ _04755_ _04798_ _04803_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__and3_2
X_13656_ clknet_leaf_64_clk _00202_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12607_ sha256cu.m_pad_pars.block_512\[15\]\[0\] _06280_ VGND VGND VPWR VPWR _06281_
+ sky130_fd_sc_hd__and2_1
X_10868_ _01976_ _04738_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__and2_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ clknet_leaf_59_clk _00133_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10799_ sha256cu.msg_scheduler.mreg_11\[26\] _04685_ _04691_ _04688_ VGND VGND VPWR
+ VPWR _00838_ sky130_fd_sc_hd__o211a_1
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12538_ sha256cu.m_pad_pars.block_512\[11\]\[1\] _06241_ VGND VGND VPWR VPWR _06243_
+ sky130_fd_sc_hd__and2_1
X_12469_ _06206_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14208_ clknet_leaf_28_clk _00754_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14139_ clknet_leaf_44_clk _00685_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06961_ _01578_ _01647_ _01613_ _01649_ _01650_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__o221a_1
X_09680_ sha256cu.iter_processing.w\[3\] _04046_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__or2_1
X_08700_ _03197_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__nor2_1
XFILLER_67_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08631_ sha256cu.m_out_digest.c_in\[14\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[14\]
+ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__o22a_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06892_ _01573_ _01577_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__and2_1
XFILLER_94_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08562_ _03155_ _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07513_ _02117_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__xnor2_2
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08493_ _03092_ _03093_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__nand2_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07444_ sha256cu.iter_processing.w\[1\] _02047_ _02046_ VGND VGND VPWR VPWR _02072_
+ sky130_fd_sc_hd__a21o_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07375_ sha256cu.counter_iteration\[0\] _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__nor2_1
X_09114_ _03567_ _03573_ _03566_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__o21ba_1
XFILLER_148_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09045_ sha256cu.m_out_digest.h_in\[14\] sha256cu.m_out_digest.d_in\[14\] VGND VGND
+ VPWR VPWR _03533_ sky130_fd_sc_hd__or2_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09947_ sha256cu.msg_scheduler.mreg_1\[12\] _04202_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__or2_1
XFILLER_104_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09878_ sha256cu.msg_scheduler.mreg_13\[24\] _04160_ VGND VGND VPWR VPWR _04164_
+ sky130_fd_sc_hd__or2_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _02230_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _05616_ _05641_ _05661_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__a21o_1
XANTENNA_303 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_325 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_314 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_347 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _05587_ _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__nor2_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_336 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_369 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ sha256cu.msg_scheduler.mreg_11\[25\] _04640_ VGND VGND VPWR VPWR _04648_
+ sky130_fd_sc_hd__or2_1
XFILLER_41_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13510_ _01975_ _06770_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__and2_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14490_ clknet_leaf_121_clk _01004_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10653_ sha256cu.msg_scheduler.mreg_10\[27\] _04601_ VGND VGND VPWR VPWR _04609_
+ sky130_fd_sc_hd__or2_1
XFILLER_41_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13441_ _04188_ _00061_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__and2b_1
X_10584_ _04529_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__buf_2
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13372_ sha256cu.m_pad_pars.block_512\[59\]\[7\] _06682_ VGND VGND VPWR VPWR _06687_
+ sky130_fd_sc_hd__and2_1
X_12323_ _06123_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12254_ _06057_ _06058_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__nand2_1
XFILLER_123_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12185_ sha256cu.msg_scheduler.mreg_1\[28\] _05992_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__xnor2_1
X_11205_ sha256cu.m_pad_pars.block_512\[22\]\[4\] _05013_ _05059_ _01970_ VGND VGND
+ VPWR VPWR _05060_ sky130_fd_sc_hd__a211o_1
XFILLER_96_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11136_ _04913_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__nor2_1
XFILLER_1_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11067_ _04747_ _04771_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__o21a_1
X_10018_ sha256cu.msg_scheduler.mreg_2\[11\] _04241_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__or2_1
XFILLER_91_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14826_ clknet_leaf_22_clk _01340_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14757_ clknet_leaf_105_clk _01271_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11969_ sha256cu.msg_scheduler.mreg_14\[3\] sha256cu.msg_scheduler.mreg_14\[1\] VGND
+ VGND VPWR VPWR _05786_ sky130_fd_sc_hd__xnor2_1
X_13708_ clknet_leaf_82_clk _00254_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[31\]
+ sky130_fd_sc_hd__dfxtp_4
X_14688_ clknet_leaf_104_clk _01202_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13639_ clknet_leaf_79_clk _00185_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07160_ _00454_ _00452_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__nor2_1
XFILLER_145_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07091_ _01663_ _01767_ _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__and3_1
XFILLER_117_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09801_ _04053_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07993_ _02604_ _02606_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__xnor2_1
X_09732_ sha256cu.iter_processing.w\[25\] _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__or2_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06944_ _01632_ _01633_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__nor2_4
XFILLER_28_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09663_ sha256cu.m_out_digest.h_in\[27\] _02369_ _02478_ sha256cu.m_out_digest.g_in\[27\]
+ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__o22a_1
XFILLER_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06875_ _01564_ _01569_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__nand2_4
XFILLER_94_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08614_ sha256cu.m_out_digest.b_in\[31\] _03177_ _03180_ sha256cu.m_out_digest.a_in\[31\]
+ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__o22a_1
X_09594_ sha256cu.m_out_digest.f_in\[31\] _04032_ _04030_ sha256cu.m_out_digest.e_in\[31\]
+ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o22a_1
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08545_ _03068_ _03071_ _03105_ _03106_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__a311o_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08476_ _03046_ _03048_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__nand2_1
XFILLER_23_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07427_ _02052_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07358_ _01993_ _01994_ _01995_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__and3b_1
XFILLER_108_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07289_ sha256cu.byte_rdy _01906_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__or2b_1
X_09028_ _03512_ _03516_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__nor2_1
XFILLER_2_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13990_ clknet_leaf_57_clk _00536_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12941_ _06458_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12872_ _06421_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_122 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ sha256cu.msg_scheduler.mreg_1\[28\] _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__xnor2_1
XANTENNA_111 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14611_ clknet_leaf_5_clk _01125_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_144 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_155 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_199 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ sha256cu.msg_scheduler.mreg_14\[24\] sha256cu.msg_scheduler.mreg_14\[17\]
+ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14542_ clknet_leaf_111_clk _01056_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_177 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11685_ _05486_ _05489_ _05485_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__a21boi_1
X_10705_ sha256cu.msg_scheduler.mreg_10\[17\] _04633_ _04638_ _04636_ VGND VGND VPWR
+ VPWR _00797_ sky130_fd_sc_hd__o211a_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ clknet_leaf_12_clk _00987_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10636_ sha256cu.msg_scheduler.mreg_9\[19\] _04594_ _04599_ _04597_ VGND VGND VPWR
+ VPWR _00767_ sky130_fd_sc_hd__o211a_1
X_13424_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10567_ sha256cu.msg_scheduler.mreg_9\[22\] _04548_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__or2_1
X_13355_ sha256cu.m_pad_pars.block_512\[58\]\[7\] _06671_ VGND VGND VPWR VPWR _06678_
+ sky130_fd_sc_hd__and2_1
X_10498_ _04414_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__clkbuf_2
X_12306_ _06107_ _06108_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__or2_1
X_13286_ sha256cu.m_pad_pars.block_512\[54\]\[6\] _06635_ VGND VGND VPWR VPWR _06642_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12237_ sha256cu.msg_scheduler.mreg_14\[14\] sha256cu.msg_scheduler.mreg_14\[12\]
+ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__xor2_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12168_ _05975_ _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__nand2_1
XFILLER_96_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12099_ _05883_ _05891_ _05910_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11119_ _04725_ _04721_ _04951_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__and3_1
Xinput6 hash[104] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14809_ clknet_leaf_117_clk _01323_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08330_ _02933_ _02895_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__a21o_1
X_08261_ _02866_ _02867_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__or2b_1
X_07212_ _01650_ _01851_ _01871_ _01874_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__o31a_1
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08192_ _02798_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__xnor2_1
X_07143_ _01705_ _01814_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__o21ai_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07074_ _00457_ _01742_ _01746_ _01754_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a31o_1
XFILLER_145_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07976_ sha256cu.K\[15\] _02581_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__nand2_1
XFILLER_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09715_ sha256cu.iter_processing.w\[18\] _04067_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__or2_1
X_06927_ _01617_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09646_ sha256cu.m_out_digest.h_in\[11\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[11\]
+ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__o22a_1
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06858_ net50 net53 net52 net55 VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__or4_1
X_06789_ net177 net181 net180 net183 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__or4_2
X_09577_ sha256cu.m_out_digest.f_in\[17\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[17\]
+ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__a22o_1
XFILLER_82_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ sha256cu.iter_processing.w\[30\] _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__xor2_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _03007_ _03008_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__and2b_1
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11470_ _01936_ _05293_ _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__and3_2
XFILLER_137_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10421_ _04396_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__buf_2
XFILLER_136_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10352_ sha256cu.msg_scheduler.mreg_5\[25\] _04434_ _04436_ _04437_ VGND VGND VPWR
+ VPWR _00645_ sky130_fd_sc_hd__o211a_1
X_13140_ _06564_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13071_ _06527_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10283_ sha256cu.msg_scheduler.mreg_5\[28\] _04387_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__or2_1
XFILLER_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12022_ _05835_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__nor2_1
X_13973_ clknet_leaf_42_clk _00519_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[27\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12924_ _06449_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__clkbuf_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _06412_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__clkbuf_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _05628_ _05629_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__nor2_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ sha256cu.m_pad_pars.block_512\[25\]\[4\] _06371_ VGND VGND VPWR VPWR _06376_
+ sky130_fd_sc_hd__and2_1
XFILLER_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11737_ _05562_ _05563_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__xnor2_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14525_ clknet_leaf_121_clk _01039_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11668_ _05473_ _05474_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__nor2_1
X_14456_ clknet_leaf_119_clk _00970_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10619_ sha256cu.msg_scheduler.mreg_10\[12\] _04588_ VGND VGND VPWR VPWR _04590_
+ sky130_fd_sc_hd__or2_1
X_14387_ clknet_leaf_47_clk _00901_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_13407_ sha256cu.m_pad_pars.m_size\[8\] sha256cu.m_pad_pars.block_512\[62\]\[0\]
+ _01923_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux2_1
X_11599_ sha256cu.flag_0_15 sha256cu.msg_scheduler.counter_iteration\[6\] sha256cu.msg_scheduler.counter_iteration\[5\]
+ _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__nor4_4
XFILLER_127_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13338_ sha256cu.m_pad_pars.block_512\[57\]\[7\] _06660_ VGND VGND VPWR VPWR _06669_
+ sky130_fd_sc_hd__and2_1
XFILLER_143_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13269_ sha256cu.m_pad_pars.block_512\[53\]\[6\] _06626_ VGND VGND VPWR VPWR _06633_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07830_ sha256cu.iter_processing.w\[12\] _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07761_ _02380_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__inv_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09500_ _03934_ _03941_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__o21a_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07692_ _02268_ _02280_ _02313_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__o21ba_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09431_ _03904_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__or2_1
XFILLER_80_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09362_ _03834_ _03839_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__or2_1
X_08313_ _02886_ _02887_ _02917_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__or3b_1
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _01526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _04881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09293_ _03734_ _03741_ _03771_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__or3_1
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_66 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ sha256cu.m_out_digest.e_in\[29\] _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__xnor2_4
XANTENNA_55 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_77 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08175_ sha256cu.m_out_digest.b_in\[21\] sha256cu.m_out_digest.a_in\[21\] _02783_
+ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_99 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07126_ _01719_ _01641_ _01696_ _01659_ _00456_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__o221a_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07057_ _01690_ _01666_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__nand2_1
XFILLER_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07959_ _02563_ _02573_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__xor2_2
X_10970_ sha256cu.m_pad_pars.block_512\[35\]\[0\] _04818_ _04822_ sha256cu.m_pad_pars.block_512\[47\]\[0\]
+ _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a221o_1
XFILLER_83_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09629_ sha256cu.m_out_digest.g_in\[29\] _04037_ _04036_ sha256cu.m_out_digest.f_in\[29\]
+ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__a22o_1
XFILLER_71_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12640_ _01912_ _05137_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__or2_2
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
X_12571_ _06251_ _04933_ _05124_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__or3_2
X_14310_ clknet_leaf_92_clk _00003_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11522_ sha256cu.m_pad_pars.block_512\[60\]\[4\] _01998_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[4\]
+ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__a22o_1
X_14241_ clknet_leaf_19_clk _00787_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11453_ _04746_ _05295_ _05277_ _01992_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__o211a_2
X_10404_ sha256cu.msg_scheduler.mreg_7\[16\] _04455_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__or2_1
X_14172_ clknet_leaf_45_clk _00718_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13123_ _06555_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__clkbuf_1
X_11384_ _05223_ _05227_ _05228_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__or3_1
X_10335_ sha256cu.msg_scheduler.mreg_5\[18\] _04421_ _04427_ _04424_ VGND VGND VPWR
+ VPWR _00638_ sky130_fd_sc_hd__o211a_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10266_ sha256cu.msg_scheduler.mreg_5\[21\] _04387_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__or2_1
XFILLER_140_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13054_ _06518_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12005_ _05775_ _05819_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__nand2_1
XFILLER_79_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10197_ sha256cu.msg_scheduler.mreg_4\[23\] _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__or2_1
XFILLER_94_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13956_ clknet_leaf_52_clk _00502_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_13887_ clknet_leaf_24_clk _00433_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12907_ sha256cu.m_pad_pars.block_512\[32\]\[5\] _06434_ VGND VGND VPWR VPWR _06440_
+ sky130_fd_sc_hd__and2_1
XFILLER_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12838_ _06403_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_41_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ sha256cu.m_pad_pars.block_512\[24\]\[4\] _06362_ VGND VGND VPWR VPWR _06367_
+ sky130_fd_sc_hd__and2_1
XFILLER_148_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14508_ clknet_leaf_12_clk _01022_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput20 hash[117] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_14439_ clknet_leaf_8_clk _00953_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput31 hash[127] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
XFILLER_30_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput42 hash[137] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 hash[157] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xinput53 hash[147] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput75 hash[167] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_116_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput97 hash[187] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xinput86 hash[177] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
X_09980_ sha256cu.msg_scheduler.mreg_1\[26\] _04215_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__or2_1
XFILLER_104_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08931_ sha256cu.m_out_digest.h_in\[10\] sha256cu.m_out_digest.d_in\[10\] VGND VGND
+ VPWR VPWR _03423_ sky130_fd_sc_hd__or2_1
X_08862_ _03343_ _03344_ _03355_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__or3_1
X_07813_ _02371_ _02393_ _02431_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__a21oi_2
XFILLER_69_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08793_ _03278_ _03276_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__or2b_1
XFILLER_57_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07744_ _02320_ _02322_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__and2b_1
X_07675_ _02294_ _02295_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__and3_1
XFILLER_53_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09414_ _03887_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__nand2_1
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
X_09345_ _03821_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__nor2_1
X_09276_ _03746_ _03747_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__nand2_1
X_08227_ _02832_ _02834_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__xor2_1
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08158_ _02761_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__nor2_1
XFILLER_107_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08089_ _02198_ _02070_ _02700_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__a21o_1
X_07109_ _01783_ _01784_ _01629_ _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__o211a_1
X_10120_ sha256cu.msg_scheduler.mreg_3\[22\] _04295_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__or2_1
X_10051_ sha256cu.msg_scheduler.mreg_1\[24\] _04260_ _04265_ _04264_ VGND VGND VPWR
+ VPWR _00516_ sky130_fd_sc_hd__o211a_1
XFILLER_88_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_99_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13810_ clknet_leaf_47_clk _00356_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14790_ clknet_leaf_116_clk _01304_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13741_ clknet_leaf_70_clk _00287_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10953_ _04779_ _04819_ _04792_ _04808_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__o22a_1
XFILLER_113_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13672_ clknet_leaf_78_clk _00218_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10884_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_23_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
X_12623_ _06270_ _05283_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__nand2_2
XFILLER_8_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12554_ _06251_ _04933_ _05295_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__or3_2
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11505_ sha256cu.data_in_padd\[26\] _01980_ _01987_ _05345_ VGND VGND VPWR VPWR _00889_
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14224_ clknet_leaf_26_clk _00770_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_12485_ sha256cu.m_pad_pars.block_512\[8\]\[0\] _06214_ VGND VGND VPWR VPWR _06215_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11436_ _04907_ _05276_ _05277_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__o211a_2
X_14155_ clknet_leaf_31_clk _00701_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11367_ sha256cu.m_pad_pars.block_512\[25\]\[5\] _05140_ _05141_ sha256cu.m_pad_pars.block_512\[29\]\[5\]
+ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__a22o_1
XFILLER_153_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14086_ clknet_leaf_37_clk _00632_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10318_ sha256cu.msg_scheduler.mreg_6\[11\] _04415_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__or2_1
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ _06546_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _06509_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__clkbuf_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ sha256cu.m_pad_pars.add_out1\[5\] sha256cu.m_pad_pars.add_out1\[4\] VGND
+ VGND VPWR VPWR _05149_ sky130_fd_sc_hd__and2_1
X_10249_ sha256cu.msg_scheduler.mreg_5\[14\] _04374_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__or2_1
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13939_ clknet_leaf_43_clk _00485_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07460_ _02082_ _02087_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__xnor2_1
X_07391_ _02019_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09130_ _03597_ _03598_ _03600_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_14_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_148_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09061_ sha256cu.K\[13\] _03515_ _03514_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__a21o_1
XFILLER_147_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08012_ _02475_ _02624_ _02625_ _02329_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__o2bb2a_1
X_09963_ _04133_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__clkbuf_2
X_08914_ sha256cu.K\[9\] _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__xor2_1
XFILLER_131_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09894_ sha256cu.msg_scheduler.mreg_12\[30\] _04167_ _04173_ _04171_ VGND VGND VPWR
+ VPWR _00445_ sky130_fd_sc_hd__o211a_1
XFILLER_57_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ sha256cu.m_out_digest.e_in\[6\] _02732_ _03339_ _03340_ _02258_ VGND VGND
+ VPWR VPWR _00229_ sky130_fd_sc_hd__a221o_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _03272_ _03273_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__nand2_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07727_ sha256cu.m_out_digest.h_in\[9\] _02347_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07658_ _02268_ _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__xor2_2
X_07589_ sha256cu.K\[5\] _02213_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09328_ _03772_ _03785_ _03806_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__and3_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09259_ sha256cu.K\[21\] _03739_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12270_ _06054_ _06056_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__a21oi_4
XFILLER_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11221_ _05024_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__and2_1
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11152_ _04771_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__nor2_2
X_10103_ _04281_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__clkbuf_2
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11083_ _04907_ _04758_ _04942_ sha256cu.m_pad_pars.block_512\[19\]\[7\] VGND VGND
+ VPWR VPWR _04943_ sky130_fd_sc_hd__o22a_1
XFILLER_1_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput210 hash[58] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10034_ sha256cu.msg_scheduler.mreg_1\[17\] _04247_ _04255_ _04250_ VGND VGND VPWR
+ VPWR _00509_ sky130_fd_sc_hd__o211a_1
Xinput254 hash[98] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput232 hash[78] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_4
Xinput243 hash[88] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
X_14911_ clknet_leaf_100_clk _01425_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[61\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput221 hash[68] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14842_ clknet_leaf_117_clk _01356_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11985_ sha256cu.msg_scheduler.mreg_1\[20\] sha256cu.msg_scheduler.mreg_1\[3\] VGND
+ VGND VPWR VPWR _05801_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14773_ clknet_leaf_3_clk _01287_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13724_ clknet_leaf_68_clk _00270_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10936_ _04785_ _04801_ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a21oi_1
X_13655_ clknet_leaf_63_clk _00201_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10867_ _04737_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__clkbuf_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _04778_ _04780_ _01912_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__a21o_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ clknet_leaf_59_clk _00132_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10798_ sha256cu.msg_scheduler.mreg_12\[26\] _04679_ VGND VGND VPWR VPWR _04691_
+ sky130_fd_sc_hd__or2_1
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12537_ _06242_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12468_ sha256cu.m_pad_pars.block_512\[7\]\[0\] _06205_ VGND VGND VPWR VPWR _06206_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14207_ clknet_leaf_45_clk _00753_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11419_ _01977_ _05125_ _05256_ _05262_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__a31o_1
X_14138_ clknet_leaf_35_clk _00684_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12399_ _01965_ _04763_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__nand2_2
XFILLER_4_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14069_ clknet_leaf_36_clk _00615_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_3_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_06960_ _01584_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__buf_2
XFILLER_140_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06891_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_4
X_08630_ sha256cu.m_out_digest.c_in\[13\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[13\]
+ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o22a_1
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08561_ _03157_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07512_ _02136_ _02138_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__xnor2_1
X_08492_ _03086_ _03091_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__or2_1
X_07443_ sha256cu.K\[2\] VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__inv_2
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09113_ _03597_ _03598_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__nor2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07374_ sha256cu.counter_iteration\[3\] sha256cu.counter_iteration\[2\] sha256cu.counter_iteration\[1\]
+ _02004_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__or4_1
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09044_ _03510_ _03511_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__nor2_1
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09946_ sha256cu.msg_scheduler.mreg_0\[11\] _04195_ _04205_ _04198_ VGND VGND VPWR
+ VPWR _00471_ sky130_fd_sc_hd__o211a_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09877_ sha256cu.msg_scheduler.mreg_12\[23\] _04153_ _04163_ _04157_ VGND VGND VPWR
+ VPWR _00438_ sky130_fd_sc_hd__o211a_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _03322_ _03323_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__nor2_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _03255_ _03257_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__xor2_1
XANTENNA_304 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_315 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_348 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_326 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _05582_ _05584_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__and2b_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_359 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_337 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10721_ sha256cu.msg_scheduler.mreg_10\[24\] _04646_ _04647_ _04636_ VGND VGND VPWR
+ VPWR _00804_ sky130_fd_sc_hd__o211a_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13440_ _06717_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__buf_2
X_10652_ sha256cu.msg_scheduler.mreg_9\[26\] _04607_ _04608_ _04597_ VGND VGND VPWR
+ VPWR _00774_ sky130_fd_sc_hd__o211a_1
XFILLER_70_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10583_ sha256cu.msg_scheduler.mreg_9\[29\] _04561_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__or2_1
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13371_ _06686_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__clkbuf_1
X_12322_ _06097_ _06100_ _06098_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__a21bo_1
X_12253_ sha256cu.msg_scheduler.mreg_9\[28\] sha256cu.msg_scheduler.mreg_0\[28\] VGND
+ VGND VPWR VPWR _06058_ sky130_fd_sc_hd__or2_1
XFILLER_107_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11204_ sha256cu.m_pad_pars.block_512\[50\]\[4\] _05008_ _04972_ sha256cu.m_pad_pars.block_512\[38\]\[4\]
+ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__a221o_1
X_12184_ sha256cu.msg_scheduler.mreg_1\[11\] sha256cu.msg_scheduler.mreg_1\[0\] VGND
+ VGND VPWR VPWR _05992_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11135_ _04701_ _04758_ _04993_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__o21a_1
XFILLER_1_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11066_ _04699_ _04924_ _04925_ sha256cu.m_pad_pars.block_512\[23\]\[7\] VGND VGND
+ VPWR VPWR _04926_ sky130_fd_sc_hd__a31o_1
X_10017_ sha256cu.msg_scheduler.mreg_1\[10\] _04234_ _04245_ _04237_ VGND VGND VPWR
+ VPWR _00502_ sky130_fd_sc_hd__o211a_1
XFILLER_92_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14825_ clknet_leaf_7_clk _01339_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14756_ clknet_leaf_106_clk _01270_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11968_ _05783_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__and2_1
X_13707_ clknet_leaf_82_clk _00253_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[30\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_60_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11899_ _05716_ _05717_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__and2_1
X_14687_ clknet_leaf_104_clk _01201_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[33\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10919_ _01943_ _04703_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__nor2_4
X_13638_ clknet_leaf_80_clk _00184_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13569_ clknet_leaf_85_clk _00115_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_07090_ _01768_ _01761_ _01751_ _01620_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__a211o_1
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07992_ _02566_ _02569_ _02605_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__o21a_1
X_09800_ sha256cu.msg_scheduler.mreg_13\[22\] _04112_ _04119_ _04117_ VGND VGND VPWR
+ VPWR _00405_ sky130_fd_sc_hd__o211a_1
X_09731_ _04053_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__buf_2
X_06943_ _01573_ _01580_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__nor2_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09662_ sha256cu.m_out_digest.h_in\[26\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[26\]
+ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__a22o_1
XFILLER_54_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06874_ sha256cu.counter_iteration\[5\] sha256cu.msg_scheduler.counter_iteration\[5\]
+ _01568_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__mux2_1
XFILLER_28_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09593_ _02515_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__buf_4
X_08613_ _02109_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__buf_4
XFILLER_55_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08544_ _03142_ _03143_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__nand2_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08475_ _03060_ _03062_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__nor2_1
XFILLER_51_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07426_ sha256cu.m_out_digest.h_in\[1\] _02054_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07357_ _01976_ _01992_ sha256cu.m_pad_pars.add_out0\[4\] VGND VGND VPWR VPWR _01995_
+ sky130_fd_sc_hd__a21o_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09027_ sha256cu.K\[13\] _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__xnor2_1
X_07288_ _01933_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09929_ sha256cu.msg_scheduler.mreg_1\[4\] _04174_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__or2_1
XFILLER_74_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12940_ sha256cu.m_pad_pars.block_512\[34\]\[4\] _06453_ VGND VGND VPWR VPWR _06458_
+ sky130_fd_sc_hd__and2_1
XFILLER_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12871_ sha256cu.m_pad_pars.block_512\[30\]\[4\] _06416_ VGND VGND VPWR VPWR _06421_
+ sky130_fd_sc_hd__and2_1
XANTENNA_123 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ sha256cu.msg_scheduler.mreg_1\[17\] sha256cu.msg_scheduler.mreg_1\[13\] VGND
+ VGND VPWR VPWR _05645_ sky130_fd_sc_hd__xnor2_1
XANTENNA_101 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ clknet_leaf_5_clk _01124_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_145 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_156 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _05577_ _05578_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__nor2_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14541_ clknet_leaf_8_clk _01055_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_178 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11684_ _05510_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__xor2_1
X_10704_ sha256cu.msg_scheduler.mreg_11\[17\] _04627_ VGND VGND VPWR VPWR _04638_
+ sky130_fd_sc_hd__or2_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ clknet_leaf_12_clk _00986_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10635_ sha256cu.msg_scheduler.mreg_10\[19\] _04588_ VGND VGND VPWR VPWR _04599_
+ sky130_fd_sc_hd__or2_1
X_13423_ sha256cu.temp_case _04177_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__nor2_4
X_13354_ _06677_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_1
X_10566_ sha256cu.msg_scheduler.mreg_8\[21\] _04554_ _04559_ _04557_ VGND VGND VPWR
+ VPWR _00737_ sky130_fd_sc_hd__o211a_1
XFILLER_115_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12305_ _06087_ _06088_ _06085_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__a21oi_1
X_10497_ sha256cu.msg_scheduler.mreg_7\[24\] _04513_ _04519_ _04516_ VGND VGND VPWR
+ VPWR _00708_ sky130_fd_sc_hd__o211a_1
XFILLER_127_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13285_ _06641_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12236_ _06040_ _06041_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__nor2_1
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12167_ _05973_ _05974_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__nand2_1
XFILLER_122_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11118_ _04913_ _04975_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__o21a_2
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12098_ _05908_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__and2b_1
Xinput7 hash[105] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
X_11049_ _04908_ _04777_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__nand2_1
XFILLER_76_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14808_ clknet_leaf_119_clk _01322_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14739_ clknet_leaf_5_clk _01253_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08260_ _02846_ _02822_ _02865_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__or3b_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08191_ sha256cu.K\[20\] _02757_ _02799_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__a21boi_2
X_07211_ _01593_ _01872_ _01873_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__a21bo_1
X_07142_ _01612_ _01703_ _01721_ _01719_ _01652_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__a221o_1
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07073_ _01749_ _01753_ _01663_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__o21a_1
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07975_ _02578_ _02580_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__or2_1
X_09714_ sha256cu.msg_scheduler.mreg_14\[17\] _04060_ _04070_ _04064_ VGND VGND VPWR
+ VPWR _00368_ sky130_fd_sc_hd__o211a_1
XFILLER_56_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06926_ _01583_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_4
X_06857_ net41 net44 net43 net47 VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__or4_2
X_09645_ sha256cu.m_out_digest.h_in\[10\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[10\]
+ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__o22a_1
XFILLER_83_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09576_ sha256cu.m_out_digest.f_in\[16\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[16\]
+ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__o22a_1
X_06788_ _01482_ _01483_ _01484_ _01485_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__or4_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _03125_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _03058_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__or2_1
X_07409_ _01913_ _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__or2_1
XFILLER_51_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10420_ sha256cu.msg_scheduler.mreg_7\[23\] _04468_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__or2_1
XFILLER_109_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08389_ _02885_ _02989_ _02992_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__o21ba_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10351_ _04396_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__buf_2
XFILLER_109_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10282_ sha256cu.msg_scheduler.mreg_4\[27\] _04393_ _04395_ _04397_ VGND VGND VPWR
+ VPWR _00615_ sky130_fd_sc_hd__o211a_1
XFILLER_117_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13070_ sha256cu.m_pad_pars.block_512\[42\]\[1\] _06525_ VGND VGND VPWR VPWR _06527_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12021_ _05807_ _05809_ _05805_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13972_ clknet_leaf_42_clk _00518_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[26\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12923_ sha256cu.m_pad_pars.block_512\[33\]\[4\] _06444_ VGND VGND VPWR VPWR _06449_
+ sky130_fd_sc_hd__and2_1
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12854_ sha256cu.m_pad_pars.block_512\[29\]\[4\] _06407_ VGND VGND VPWR VPWR _06412_
+ sky130_fd_sc_hd__and2_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _05626_ _05627_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__and2_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12785_ _06375_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__clkbuf_1
X_11736_ _05538_ _05541_ _05537_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__a21oi_2
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14524_ clknet_leaf_126_clk _01038_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ _05494_ _05496_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__xnor2_1
X_14455_ clknet_leaf_120_clk _00969_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10618_ sha256cu.msg_scheduler.mreg_9\[11\] _04581_ _04589_ _04584_ VGND VGND VPWR
+ VPWR _00759_ sky130_fd_sc_hd__o211a_1
X_14386_ clknet_leaf_47_clk _00900_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_13406_ _06704_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__clkbuf_1
X_11598_ sha256cu.msg_scheduler.counter_iteration\[4\] _01565_ _04716_ VGND VGND VPWR
+ VPWR _05431_ sky130_fd_sc_hd__a21o_1
X_10549_ sha256cu.msg_scheduler.mreg_9\[14\] _04548_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__or2_1
XFILLER_6_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13337_ _06668_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13268_ _06632_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12219_ _06024_ _06025_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__or2_1
X_13199_ sha256cu.m_pad_pars.block_512\[49\]\[5\] _06590_ VGND VGND VPWR VPWR _06596_
+ sky130_fd_sc_hd__and2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07760_ sha256cu.m_out_digest.e_in\[21\] _02379_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__xnor2_2
XFILLER_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07691_ _02277_ _02279_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__nor2_1
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09430_ _03902_ _03903_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__and2_1
XFILLER_80_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09361_ _03725_ _03780_ _03835_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__o31a_1
X_09292_ _03734_ _03741_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__o21ai_1
X_08312_ _02886_ _02887_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__o21ba_1
X_08243_ sha256cu.m_out_digest.e_in\[16\] sha256cu.m_out_digest.e_in\[2\] VGND VGND
+ VPWR VPWR _02850_ sky130_fd_sc_hd__xnor2_4
XANTENNA_12 _01551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _05342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_67 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ sha256cu.m_out_digest.b_in\[21\] sha256cu.m_out_digest.a_in\[21\] sha256cu.m_out_digest.c_in\[21\]
+ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__a21o_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07125_ _01761_ _01795_ _01796_ _01798_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__o32a_1
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07056_ _01642_ _01639_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__nor2_1
XFILLER_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07958_ _02570_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__xnor2_2
XFILLER_75_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07889_ _02461_ _02459_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__and2b_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06909_ _01592_ _00453_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__nor2_2
XFILLER_83_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09628_ sha256cu.m_out_digest.g_in\[28\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[28\]
+ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__o22a_1
XFILLER_71_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09559_ _02109_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__buf_4
XFILLER_24_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12570_ _06260_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11521_ sha256cu.m_pad_pars.block_512\[20\]\[4\] _05294_ _05285_ sha256cu.m_pad_pars.block_512\[16\]\[4\]
+ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a22o_1
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14240_ clknet_leaf_19_clk _00786_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11452_ _04701_ _05248_ _04751_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__o21a_1
X_10403_ sha256cu.msg_scheduler.mreg_6\[15\] _04461_ _04466_ _04464_ VGND VGND VPWR
+ VPWR _00667_ sky130_fd_sc_hd__o211a_1
X_14171_ clknet_leaf_45_clk _00717_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11383_ sha256cu.m_pad_pars.block_512\[41\]\[6\] _05132_ _05147_ sha256cu.m_pad_pars.block_512\[33\]\[6\]
+ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__a22o_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10334_ sha256cu.msg_scheduler.mreg_6\[18\] _04415_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__or2_1
X_13122_ sha256cu.m_pad_pars.block_512\[45\]\[1\] _06553_ VGND VGND VPWR VPWR _06555_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10265_ _04281_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__clkbuf_2
XFILLER_140_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13053_ sha256cu.m_pad_pars.block_512\[41\]\[1\] _06516_ VGND VGND VPWR VPWR _06518_
+ sky130_fd_sc_hd__and2_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10196_ _04281_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__clkbuf_2
X_12004_ _05794_ _05813_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__and2_1
XFILLER_79_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13955_ clknet_leaf_52_clk _00501_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_81_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13886_ clknet_leaf_24_clk _00432_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12906_ _06439_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__clkbuf_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ sha256cu.m_pad_pars.block_512\[28\]\[4\] _06398_ VGND VGND VPWR VPWR _06403_
+ sky130_fd_sc_hd__and2_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _06366_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11719_ _05521_ _05525_ _05545_ _05432_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__a31o_1
X_14507_ clknet_leaf_8_clk _01021_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12699_ _06329_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_1
Xinput10 hash[108] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 hash[118] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
X_14438_ clknet_leaf_103_clk _00952_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput43 hash[138] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput54 hash[148] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xinput32 hash[128] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput76 hash[168] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
Xinput98 hash[188] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
X_14369_ clknet_leaf_77_clk _00883_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput87 hash[178] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput65 hash[158] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08930_ _03410_ _03411_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__nand2_1
XFILLER_130_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08861_ _03343_ _03344_ _03355_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07812_ _02392_ _02390_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__and2b_1
XFILLER_69_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08792_ _03289_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__inv_1
X_07743_ _02362_ _02363_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__nand2_1
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07674_ sha256cu.m_out_digest.g_in\[8\] sha256cu.m_out_digest.f_in\[8\] sha256cu.m_out_digest.e_in\[8\]
+ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__mux2_1
XFILLER_93_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09413_ _03860_ _03861_ _03888_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a21bo_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09344_ sha256cu.iter_processing.w\[24\] _02903_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__and2_1
XFILLER_40_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09275_ _02332_ _03754_ _03755_ _03366_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__o211a_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08226_ _02772_ _02791_ _02833_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__o21ai_1
X_08157_ _02627_ _02763_ _02766_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__o21a_1
XFILLER_147_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07108_ _01657_ _01580_ _01653_ _01734_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__a31o_1
XFILLER_106_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08088_ _02695_ _02698_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__o21a_1
XFILLER_115_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07039_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__inv_2
X_10050_ sha256cu.msg_scheduler.mreg_2\[24\] _04254_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__or2_1
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13740_ clknet_leaf_70_clk _00286_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10952_ sha256cu.m_pad_pars.add_512_block\[6\] _04791_ VGND VGND VPWR VPWR _04819_
+ sky130_fd_sc_hd__or2_2
XFILLER_83_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13671_ clknet_leaf_80_clk _00217_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10883_ _04748_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__or2_1
X_12622_ _01966_ _04938_ _06288_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a21oi_1
X_12553_ _01911_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__buf_4
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11504_ _05337_ _05339_ _05344_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__or3_2
XFILLER_12_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14223_ clknet_leaf_26_clk _00769_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[21\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12484_ _01965_ _05317_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__nand2_2
X_11435_ sha256cu.m_pad_pars.add_out0\[2\] sha256cu.m_pad_pars.add_out0\[3\] VGND
+ VGND VPWR VPWR _05278_ sky130_fd_sc_hd__nor2b_2
XFILLER_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14154_ clknet_leaf_31_clk _00700_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11366_ sha256cu.m_pad_pars.block_512\[13\]\[5\] _05128_ _05132_ sha256cu.m_pad_pars.block_512\[41\]\[5\]
+ _05211_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__a221o_1
XFILLER_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14085_ clknet_leaf_37_clk _00631_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10317_ sha256cu.msg_scheduler.mreg_5\[10\] _04407_ _04417_ _04410_ VGND VGND VPWR
+ VPWR _00630_ sky130_fd_sc_hd__o211a_1
XFILLER_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13105_ sha256cu.m_pad_pars.block_512\[44\]\[1\] _06544_ VGND VGND VPWR VPWR _06546_
+ sky130_fd_sc_hd__and2_1
X_11297_ sha256cu.m_pad_pars.block_512\[9\]\[0\] _05144_ _05147_ sha256cu.m_pad_pars.block_512\[33\]\[0\]
+ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__a22o_1
X_10248_ sha256cu.msg_scheduler.mreg_4\[13\] _04367_ _04377_ _04370_ VGND VGND VPWR
+ VPWR _00601_ sky130_fd_sc_hd__o211a_1
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ sha256cu.m_pad_pars.block_512\[40\]\[1\] _06507_ VGND VGND VPWR VPWR _06509_
+ sky130_fd_sc_hd__and2_1
XFILLER_140_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10179_ sha256cu.msg_scheduler.mreg_3\[15\] _04328_ _04338_ _04331_ VGND VGND VPWR
+ VPWR _00571_ sky130_fd_sc_hd__o211a_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13938_ clknet_leaf_50_clk _00484_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13869_ clknet_leaf_20_clk _00415_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07390_ sha256cu.m_out_digest.g_in\[0\] sha256cu.m_out_digest.f_in\[0\] sha256cu.m_out_digest.e_in\[0\]
+ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__mux2_1
XFILLER_148_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09060_ _03546_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__and2_1
XFILLER_148_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08011_ _02402_ _02471_ _02546_ _02622_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__nand4_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09962_ sha256cu.msg_scheduler.mreg_0\[18\] _04208_ _04214_ _04211_ VGND VGND VPWR
+ VPWR _00478_ sky130_fd_sc_hd__o211a_1
XFILLER_89_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08913_ _03404_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__nand2_1
XFILLER_131_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09893_ sha256cu.msg_scheduler.mreg_13\[30\] _04160_ VGND VGND VPWR VPWR _04173_
+ sky130_fd_sc_hd__or2_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _03315_ _03338_ _02732_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ sha256cu.iter_processing.w\[4\] _02153_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__nand2_1
XFILLER_57_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07726_ sha256cu.m_out_digest.a_in\[31\] _02346_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__xnor2_4
XFILLER_73_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07657_ _02277_ _02279_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__xnor2_2
XFILLER_81_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07588_ _02210_ _02212_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__xor2_1
XFILLER_43_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09327_ _03804_ _03805_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__xnor2_1
X_09258_ _03737_ _03738_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__nor2_1
XFILLER_135_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09189_ sha256cu.m_out_digest.h_in\[19\] sha256cu.m_out_digest.d_in\[19\] VGND VGND
+ VPWR VPWR _03672_ sky130_fd_sc_hd__nand2_1
X_08209_ sha256cu.m_out_digest.b_in\[22\] _02026_ sha256cu.m_out_digest.c_in\[22\]
+ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__a21o_1
XFILLER_153_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11220_ sha256cu.m_pad_pars.block_512\[62\]\[6\] _04984_ _04982_ sha256cu.m_pad_pars.block_512\[58\]\[6\]
+ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__a22o_1
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11151_ _04699_ _04925_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__nand2_1
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10102_ sha256cu.msg_scheduler.mreg_2\[14\] _04288_ _04294_ _04291_ VGND VGND VPWR
+ VPWR _00538_ sky130_fd_sc_hd__o211a_1
Xinput211 hash[59] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
Xinput200 hash[49] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11082_ _04761_ _04807_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__nor2_1
XFILLER_1_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput222 hash[69] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
X_10033_ sha256cu.msg_scheduler.mreg_2\[17\] _04254_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__or2_1
Xinput233 hash[79] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14910_ clknet_leaf_117_clk _01424_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput244 hash[89] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_2
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput255 hash[99] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_2
X_14841_ clknet_leaf_118_clk _01355_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11984_ _05798_ _05799_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__nand2_1
XFILLER_91_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14772_ clknet_leaf_3_clk _01286_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13723_ clknet_leaf_67_clk _00269_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10935_ _04751_ _04794_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__nor2_1
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13654_ clknet_leaf_63_clk _00200_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10866_ sha256cu.m_pad_pars.add_out3\[3\] sha256cu.m_pad_pars.add_out3\[2\] _04736_
+ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__and3_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12605_ _06279_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13585_ clknet_leaf_51_clk _00131_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10797_ sha256cu.msg_scheduler.mreg_11\[25\] _04685_ _04690_ _04688_ VGND VGND VPWR
+ VPWR _00837_ sky130_fd_sc_hd__o211a_1
XFILLER_40_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12536_ sha256cu.m_pad_pars.block_512\[11\]\[0\] _06241_ VGND VGND VPWR VPWR _06242_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12467_ _01912_ _04773_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__or2_2
XFILLER_125_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14206_ clknet_leaf_45_clk _00752_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11418_ _01977_ _05127_ _05258_ _05261_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__a31o_1
X_14137_ clknet_leaf_34_clk _00683_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12398_ _01966_ _05119_ _06168_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11349_ sha256cu.m_pad_pars.block_512\[53\]\[3\] _05161_ _05165_ sha256cu.m_pad_pars.block_512\[37\]\[3\]
+ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__a221o_1
XFILLER_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14068_ clknet_leaf_38_clk _00614_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06890_ _01583_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_4
X_13019_ sha256cu.m_pad_pars.block_512\[39\]\[1\] _06498_ VGND VGND VPWR VPWR _06500_
+ sky130_fd_sc_hd__and2_1
XFILLER_67_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08560_ sha256cu.iter_processing.w\[31\] _03158_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__xnor2_1
X_07511_ _02079_ _02091_ _02137_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__o21ba_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08491_ _03086_ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__nand2_1
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07442_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__buf_4
XFILLER_22_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07373_ sha256cu.iter_processing.temp_case _02006_ _02007_ sha256cu.iter_processing.temp_if
+ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__a31o_1
XFILLER_148_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09112_ _03592_ _03596_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__and2_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09043_ _03522_ _03523_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__nand2_1
XFILLER_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09945_ sha256cu.msg_scheduler.mreg_1\[11\] _04202_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__or2_1
XFILLER_98_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09876_ sha256cu.msg_scheduler.mreg_13\[23\] _04160_ VGND VGND VPWR VPWR _04163_
+ sky130_fd_sc_hd__or2_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ sha256cu.m_out_digest.h_in\[6\] sha256cu.m_out_digest.d_in\[6\] VGND VGND
+ VPWR VPWR _03323_ sky130_fd_sc_hd__and2_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _03221_ _03235_ _03256_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__a21boi_1
XANTENNA_316 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_305 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_349 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_327 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _02323_ _02329_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__or2_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ sha256cu.m_out_digest.d_in\[30\] _03189_ _03192_ sha256cu.m_out_digest.c_in\[30\]
+ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__a22o_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_338 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ sha256cu.msg_scheduler.mreg_11\[24\] _04640_ VGND VGND VPWR VPWR _04647_
+ sky130_fd_sc_hd__or2_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10651_ sha256cu.msg_scheduler.mreg_10\[26\] _04601_ VGND VGND VPWR VPWR _04608_
+ sky130_fd_sc_hd__or2_1
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10582_ sha256cu.msg_scheduler.mreg_8\[28\] _04567_ _04568_ _04557_ VGND VGND VPWR
+ VPWR _00744_ sky130_fd_sc_hd__o211a_1
X_13370_ sha256cu.m_pad_pars.block_512\[59\]\[6\] _06682_ VGND VGND VPWR VPWR _06686_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12321_ _06120_ _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__xnor2_1
X_12252_ sha256cu.msg_scheduler.mreg_9\[28\] sha256cu.msg_scheduler.mreg_0\[28\] VGND
+ VGND VPWR VPWR _06057_ sky130_fd_sc_hd__nand2_1
XFILLER_123_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11203_ sha256cu.m_pad_pars.block_512\[34\]\[4\] _04996_ _04981_ sha256cu.m_pad_pars.block_512\[54\]\[4\]
+ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__a22o_1
X_12183_ _05989_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__nand2_1
XFILLER_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11134_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__buf_2
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11065_ _04701_ _04744_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__nor2_1
X_10016_ sha256cu.msg_scheduler.mreg_2\[10\] _04241_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__or2_1
XFILLER_135_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14824_ clknet_leaf_9_clk _01338_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11967_ _05781_ _05782_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__nand2_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14755_ clknet_leaf_103_clk _01269_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13706_ clknet_leaf_82_clk _00252_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[29\]
+ sky130_fd_sc_hd__dfxtp_4
X_10918_ _04749_ _04752_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__nor2_2
X_11898_ _05716_ _05717_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__nor2_1
XFILLER_71_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14686_ clknet_leaf_115_clk _01200_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10849_ _04724_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
X_13637_ clknet_leaf_81_clk _00183_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13568_ clknet_leaf_69_clk _00114_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12519_ sha256cu.m_pad_pars.block_512\[10\]\[0\] _06232_ VGND VGND VPWR VPWR _06233_
+ sky130_fd_sc_hd__and2_1
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13499_ sha256cu.K\[25\] _06716_ _06717_ _06763_ _06737_ VGND VGND VPWR VPWR _01466_
+ sky130_fd_sc_hd__o221a_1
XFILLER_141_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07991_ sha256cu.m_out_digest.h_in\[15\] _02568_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__nand2_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09730_ sha256cu.msg_scheduler.mreg_14\[24\] _04073_ _04079_ _04077_ VGND VGND VPWR
+ VPWR _00375_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_06942_ _01573_ _01577_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__nor2_4
XFILLER_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09661_ sha256cu.m_out_digest.h_in\[25\] _02369_ _02478_ sha256cu.m_out_digest.g_in\[25\]
+ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__o22a_1
X_06873_ sha256cu.msg_scheduler.temp_case _01567_ sha256cu.iter_processing.padding_done
+ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__o21a_2
XFILLER_131_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08612_ sha256cu.m_out_digest.b_in\[30\] _03179_ _03178_ _02304_ VGND VGND VPWR VPWR
+ _00157_ sky130_fd_sc_hd__a22o_1
X_09592_ sha256cu.m_out_digest.f_in\[30\] _04029_ _04031_ sha256cu.m_out_digest.e_in\[30\]
+ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__a22o_1
XFILLER_55_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08543_ _03101_ _03112_ _03141_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__or3b_1
XFILLER_54_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08474_ sha256cu.K\[29\] VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__clkinv_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07425_ sha256cu.m_out_digest.a_in\[23\] _02053_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__xnor2_2
XFILLER_51_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07356_ _01964_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__buf_4
XFILLER_149_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07287_ sha256cu.m_pad_pars.m_size\[7\] sha256cu.m_pad_pars.block_512\[63\]\[7\]
+ _01923_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__mux2_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09026_ _03513_ _03514_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__nor2_1
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09928_ _04166_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09859_ _04044_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__buf_2
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12870_ _06420_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_124 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _05642_ _05643_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__nand2_1
XANTENNA_102 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_146 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14540_ clknet_leaf_11_clk _01054_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_135 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11752_ _05575_ _05576_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__and2_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_168 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11683_ sha256cu.msg_scheduler.mreg_1\[22\] _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__xnor2_2
X_10703_ sha256cu.msg_scheduler.mreg_10\[16\] _04633_ _04637_ _04636_ VGND VGND VPWR
+ VPWR _00796_ sky130_fd_sc_hd__o211a_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ clknet_leaf_13_clk _00985_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10634_ sha256cu.msg_scheduler.mreg_9\[18\] _04594_ _04598_ _04597_ VGND VGND VPWR
+ VPWR _00766_ sky130_fd_sc_hd__o211a_1
X_13422_ _06712_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_1
X_13353_ sha256cu.m_pad_pars.block_512\[58\]\[6\] _06671_ VGND VGND VPWR VPWR _06677_
+ sky130_fd_sc_hd__and2_1
XFILLER_139_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10565_ sha256cu.msg_scheduler.mreg_9\[21\] _04548_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__or2_1
X_12304_ _06105_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__nand2_1
X_10496_ sha256cu.msg_scheduler.mreg_8\[24\] _04507_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__or2_1
X_13284_ sha256cu.m_pad_pars.block_512\[54\]\[5\] _06635_ VGND VGND VPWR VPWR _06641_
+ sky130_fd_sc_hd__and2_1
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12235_ _06038_ _06039_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__and2_1
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12166_ _05973_ _05974_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__or2_1
XFILLER_69_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11117_ _04720_ _04966_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__nor2_1
X_12097_ _05874_ _05879_ _05907_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__a21o_1
Xinput8 hash[106] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
X_11048_ _04704_ _04744_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__nor2_4
XFILLER_76_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14807_ clknet_leaf_119_clk _01321_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[48\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12999_ _06270_ _04971_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__nand2_2
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14738_ clknet_leaf_9_clk _01252_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14669_ clknet_leaf_12_clk _01183_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_08190_ _02756_ _02735_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__or2b_1
X_07210_ _01622_ _01639_ _01658_ _01584_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__o31a_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07141_ _01594_ _01666_ _00455_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__a21oi_1
X_07072_ _01625_ _01620_ _01653_ _01635_ _01752_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__a41o_1
XFILLER_126_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07974_ _02084_ _02220_ _02587_ _02588_ _02258_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__a221o_1
XFILLER_102_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09713_ sha256cu.iter_processing.w\[17\] _04067_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__or2_1
X_06925_ _01615_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__inv_2
X_09644_ sha256cu.m_out_digest.h_in\[9\] _04037_ _04040_ sha256cu.m_out_digest.g_in\[9\]
+ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__a22o_1
XFILLER_110_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06856_ net46 net49 net48 net51 VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__or4_4
XFILLER_83_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06787_ net204 net207 net206 net209 VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__or4_2
X_09575_ sha256cu.m_out_digest.f_in\[15\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[15\]
+ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__a22o_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ sha256cu.m_out_digest.g_in\[30\] sha256cu.m_out_digest.f_in\[30\] sha256cu.m_out_digest.e_in\[30\]
+ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__mux2_2
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08457_ _03040_ _03011_ _03057_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__and3_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07408_ _02017_ _02035_ _02036_ _02037_ sha256cu.m_out_digest.a_in\[0\] VGND VGND
+ VPWR VPWR _02038_ sky130_fd_sc_hd__a32o_1
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08388_ _02918_ _02990_ _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__o21a_1
XFILLER_137_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07339_ _01980_ _01968_ sha256cu.m_pad_pars.add_out1\[4\] VGND VGND VPWR VPWR _01981_
+ sky130_fd_sc_hd__or3b_1
X_10350_ sha256cu.msg_scheduler.mreg_6\[25\] _04428_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__or2_1
XFILLER_152_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10281_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__buf_2
X_09009_ _03443_ _03471_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__nand2_1
XFILLER_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _05833_ _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__nand2_1
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13971_ clknet_leaf_42_clk _00517_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[25\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12922_ _06448_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _06411_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _05626_ _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__nor2_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ sha256cu.m_pad_pars.block_512\[25\]\[3\] _06371_ VGND VGND VPWR VPWR _06375_
+ sky130_fd_sc_hd__and2_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _05560_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__nand2_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14523_ clknet_leaf_125_clk _01037_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ clknet_leaf_112_clk _00968_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11666_ sha256cu.msg_scheduler.mreg_14\[22\] _05495_ VGND VGND VPWR VPWR _05496_
+ sky130_fd_sc_hd__xnor2_1
X_13405_ sha256cu.m_pad_pars.block_512\[61\]\[7\] _01928_ VGND VGND VPWR VPWR _06704_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10617_ sha256cu.msg_scheduler.mreg_10\[11\] _04588_ VGND VGND VPWR VPWR _04589_
+ sky130_fd_sc_hd__or2_1
X_11597_ _04580_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__clkbuf_4
X_14385_ clknet_leaf_47_clk _00899_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_143_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10548_ sha256cu.msg_scheduler.mreg_8\[13\] _04540_ _04549_ _04543_ VGND VGND VPWR
+ VPWR _00729_ sky130_fd_sc_hd__o211a_1
X_13336_ sha256cu.m_pad_pars.block_512\[57\]\[6\] _06660_ VGND VGND VPWR VPWR _06668_
+ sky130_fd_sc_hd__and2_1
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13267_ sha256cu.m_pad_pars.block_512\[53\]\[5\] _06626_ VGND VGND VPWR VPWR _06632_
+ sky130_fd_sc_hd__and2_1
X_10479_ sha256cu.msg_scheduler.mreg_7\[16\] _04500_ _04509_ _04503_ VGND VGND VPWR
+ VPWR _00700_ sky130_fd_sc_hd__o211a_1
X_12218_ _05996_ _06000_ _06023_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__and3_1
X_13198_ _06595_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12149_ sha256cu.data_in_padd\[23\] _05447_ _04692_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__a21o_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07690_ _02300_ _02311_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__xor2_2
XFILLER_65_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09360_ _03777_ _03807_ _03835_ _03836_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__o221a_1
X_09291_ _03769_ _03770_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__nor2_1
X_08311_ _02888_ _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__xnor2_1
XANTENNA_13 _01551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08242_ sha256cu.m_out_digest.h_in\[23\] _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__xnor2_1
XANTENNA_24 sha256cu.iter_processing.w\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08173_ _02778_ _02781_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__xor2_1
XFILLER_137_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07124_ _01657_ _01627_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__nor2_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07055_ _01657_ _01653_ _01611_ _01642_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o31a_1
XFILLER_88_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07957_ _02526_ _02529_ _02571_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__o21a_1
X_06908_ _01600_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkinv_2
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07888_ _02485_ _02504_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09627_ sha256cu.m_out_digest.g_in\[27\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[27\]
+ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__o22a_1
XFILLER_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06839_ _01533_ _01534_ _01535_ _01536_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__or4_2
X_09558_ sha256cu.m_out_digest.f_in\[2\] _03191_ _03190_ sha256cu.m_out_digest.e_in\[2\]
+ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__o22a_1
X_08509_ _03068_ _03071_ _03108_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09489_ _03045_ _03930_ _03929_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__a21boi_1
X_11520_ sha256cu.m_pad_pars.block_512\[12\]\[4\] _05299_ _05304_ sha256cu.m_pad_pars.block_512\[36\]\[4\]
+ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__a221o_1
XFILLER_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11451_ _04907_ _05292_ _05293_ _05277_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__o211a_2
X_10402_ sha256cu.msg_scheduler.mreg_7\[15\] _04455_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__or2_1
X_14170_ clknet_leaf_35_clk _00716_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11382_ sha256cu.m_pad_pars.block_512\[49\]\[6\] _05151_ _05158_ sha256cu.m_pad_pars.block_512\[21\]\[6\]
+ _05226_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__a221o_1
X_10333_ sha256cu.msg_scheduler.mreg_5\[17\] _04421_ _04426_ _04424_ VGND VGND VPWR
+ VPWR _00637_ sky130_fd_sc_hd__o211a_1
X_13121_ _06554_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10264_ sha256cu.msg_scheduler.mreg_4\[20\] _04380_ _04386_ _04383_ VGND VGND VPWR
+ VPWR _00608_ sky130_fd_sc_hd__o211a_1
XFILLER_112_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13052_ _06517_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__clkbuf_1
X_10195_ sha256cu.msg_scheduler.mreg_3\[22\] _04341_ _04347_ _04344_ VGND VGND VPWR
+ VPWR _00578_ sky130_fd_sc_hd__o211a_1
X_12003_ _05792_ _05812_ _05811_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__a21o_1
XFILLER_66_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13954_ clknet_leaf_54_clk _00500_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13885_ clknet_leaf_24_clk _00431_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12905_ sha256cu.m_pad_pars.block_512\[32\]\[4\] _06434_ VGND VGND VPWR VPWR _06439_
+ sky130_fd_sc_hd__and2_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ _06402_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__clkbuf_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14506_ clknet_leaf_16_clk _01020_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ sha256cu.m_pad_pars.block_512\[24\]\[3\] _06362_ VGND VGND VPWR VPWR _06366_
+ sky130_fd_sc_hd__and2_1
X_11718_ _05521_ _05525_ _05545_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__a21oi_1
X_12698_ sha256cu.m_pad_pars.block_512\[20\]\[3\] _06325_ VGND VGND VPWR VPWR _06329_
+ sky130_fd_sc_hd__and2_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11649_ _05466_ _05467_ _05478_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__nand3_1
Xinput11 hash[109] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 hash[119] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
X_14437_ clknet_leaf_97_clk _00951_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput44 hash[139] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput33 hash[129] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
X_14368_ clknet_leaf_77_clk _00882_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput55 hash[149] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput88 hash[179] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput77 hash[169] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 hash[159] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
X_13319_ sha256cu.m_pad_pars.block_512\[56\]\[6\] _01924_ VGND VGND VPWR VPWR _06659_
+ sky130_fd_sc_hd__and2_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14299_ clknet_leaf_97_clk _00011_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__dfxtp_1
Xinput99 hash[189] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08860_ _03348_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__xor2_1
XFILLER_130_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07811_ _02410_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__xnor2_2
X_08791_ _03261_ _02440_ _03286_ _03287_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__o221a_1
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07742_ _02334_ _02361_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__or2_1
XFILLER_26_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07673_ sha256cu.m_out_digest.b_in\[8\] sha256cu.m_out_digest.a_in\[8\] sha256cu.m_out_digest.c_in\[8\]
+ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__a21o_1
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09412_ _03859_ _03858_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__or2b_1
XFILLER_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09343_ sha256cu.iter_processing.w\[24\] _02903_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__nor2_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09274_ sha256cu.m_out_digest.e_in\[21\] _02439_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__or2_1
XFILLER_21_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08225_ _02788_ _02790_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__or2_1
XFILLER_32_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08156_ _02729_ _02764_ _02762_ _02697_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__a221oi_4
XFILLER_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07107_ _01603_ _01594_ _01666_ _01617_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__a31o_1
XFILLER_146_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08087_ _02695_ _02698_ _02108_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__a21oi_1
XFILLER_121_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07038_ _01667_ _01590_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__nor2_2
XFILLER_130_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08989_ _02450_ _03478_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10951_ sha256cu.m_pad_pars.add_out3\[3\] sha256cu.m_pad_pars.add_out3\[2\] _04814_
+ _04817_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__nor4_4
XFILLER_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ clknet_leaf_80_clk _00216_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12621_ _03288_ sha256cu.m_pad_pars.block_512\[15\]\[7\] VGND VGND VPWR VPWR _06288_
+ sky130_fd_sc_hd__nor2_1
XFILLER_44_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10882_ sha256cu.m_pad_pars.add_512_block\[2\] sha256cu.m_pad_pars.add_512_block\[3\]
+ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__or2b_1
XFILLER_43_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12552_ _06250_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11503_ sha256cu.m_pad_pars.block_512\[0\]\[2\] _05314_ _05340_ _05343_ VGND VGND
+ VPWR VPWR _05344_ sky130_fd_sc_hd__a211o_1
XFILLER_12_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12483_ _06213_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14222_ clknet_leaf_26_clk _00768_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[20\]
+ sky130_fd_sc_hd__dfxtp_2
X_11434_ sha256cu.m_pad_pars.add_out0\[5\] sha256cu.m_pad_pars.add_out0\[4\] VGND
+ VGND VPWR VPWR _05277_ sky130_fd_sc_hd__nor2b_2
XFILLER_153_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14153_ clknet_leaf_31_clk _00699_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11365_ sha256cu.m_pad_pars.block_512\[45\]\[5\] _05126_ VGND VGND VPWR VPWR _05211_
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_100_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_16
X_14084_ clknet_leaf_37_clk _00630_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10316_ sha256cu.msg_scheduler.mreg_6\[10\] _04415_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__or2_1
XFILLER_113_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13104_ _06545_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__clkbuf_1
X_11296_ _05125_ _05134_ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__and3_2
X_10247_ sha256cu.msg_scheduler.mreg_5\[13\] _04374_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__or2_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _06508_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__clkbuf_1
X_10178_ sha256cu.msg_scheduler.mreg_4\[15\] _04335_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__or2_1
XFILLER_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13937_ clknet_leaf_53_clk _00483_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13868_ clknet_leaf_18_clk _00414_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13799_ clknet_leaf_83_clk _00345_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12819_ _06393_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08010_ _02546_ _02622_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__and2_1
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09961_ sha256cu.msg_scheduler.mreg_1\[18\] _04202_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__or2_1
XFILLER_103_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08912_ sha256cu.iter_processing.w\[9\] _02338_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__nand2_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09892_ sha256cu.msg_scheduler.mreg_12\[29\] _04167_ _04172_ _04171_ VGND VGND VPWR
+ VPWR _00444_ sky130_fd_sc_hd__o211a_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _03315_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__or2_1
XFILLER_84_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ sha256cu.iter_processing.w\[4\] _02153_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__or2_1
XFILLER_85_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07725_ _02026_ sha256cu.m_out_digest.a_in\[11\] VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__xnor2_2
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07656_ _02231_ _02236_ _02278_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__o21a_1
XFILLER_81_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07587_ _02150_ _02173_ _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09326_ sha256cu.K\[22\] _03767_ _03766_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__a21o_1
X_09257_ sha256cu.iter_processing.w\[21\] _02785_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__and2_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08208_ _02812_ _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09188_ sha256cu.m_out_digest.h_in\[19\] sha256cu.m_out_digest.d_in\[19\] VGND VGND
+ VPWR VPWR _03671_ sky130_fd_sc_hd__or2_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08139_ sha256cu.m_out_digest.h_in\[19\] _02715_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__nand2_1
XFILLER_150_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11150_ _04747_ _04975_ _04727_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__o21a_2
XFILLER_1_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10101_ sha256cu.msg_scheduler.mreg_3\[14\] _04282_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__or2_1
XFILLER_122_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11081_ _04764_ _04766_ _04935_ _04940_ _01970_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__a311o_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput201 hash[4] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_2
Xinput223 hash[6] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
Xinput234 hash[7] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
X_10032_ _04133_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__clkbuf_2
XFILLER_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput212 hash[5] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput245 hash[8] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_4
Xinput256 hash[9] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14840_ clknet_leaf_119_clk _01354_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14771_ clknet_leaf_3_clk _01285_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11983_ sha256cu.msg_scheduler.mreg_9\[17\] sha256cu.msg_scheduler.mreg_0\[17\] VGND
+ VGND VPWR VPWR _05799_ sky130_fd_sc_hd__nand2_1
X_13722_ clknet_leaf_67_clk _00268_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10934_ _04704_ _04791_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nor2_4
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13653_ clknet_leaf_61_clk _00199_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10865_ sha256cu.m_pad_pars.add_out3\[5\] sha256cu.m_pad_pars.add_out3\[4\] VGND
+ VGND VPWR VPWR _04736_ sky130_fd_sc_hd__and2_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ clknet_leaf_51_clk _00130_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12604_ sha256cu.m_pad_pars.block_512\[14\]\[7\] _05097_ _06249_ VGND VGND VPWR VPWR
+ _06279_ sky130_fd_sc_hd__mux2_1
XFILLER_31_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10796_ sha256cu.msg_scheduler.mreg_12\[25\] _04679_ VGND VGND VPWR VPWR _04690_
+ sky130_fd_sc_hd__or2_1
X_12535_ _01965_ _04789_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__nand2_2
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12466_ _06204_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14205_ clknet_leaf_45_clk _00751_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12397_ _03288_ sha256cu.m_pad_pars.block_512\[2\]\[7\] VGND VGND VPWR VPWR _06168_
+ sky130_fd_sc_hd__nor2_1
X_11417_ _05127_ _05139_ _05260_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__and3_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14136_ clknet_leaf_34_clk _00682_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11348_ sha256cu.m_pad_pars.block_512\[5\]\[3\] _05160_ _05195_ _05024_ VGND VGND
+ VPWR VPWR _05196_ sky130_fd_sc_hd__a22o_1
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14067_ clknet_leaf_38_clk _00613_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11279_ _04702_ _04960_ _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__o21a_1
XFILLER_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13018_ _06499_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07510_ _02088_ _02090_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nor2_1
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08490_ sha256cu.iter_processing.w\[29\] _03090_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__xor2_1
X_07441_ _02065_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__buf_6
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07372_ _01964_ sha256cu.iter_processing.padding_done VGND VGND VPWR VPWR _02007_
+ sky130_fd_sc_hd__and2_1
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09111_ _03592_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__nor2_1
XFILLER_31_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09042_ _03528_ _03529_ _03530_ _03366_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__o211a_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09944_ sha256cu.msg_scheduler.mreg_0\[10\] _04195_ _04204_ _04198_ VGND VGND VPWR
+ VPWR _00470_ sky130_fd_sc_hd__o211a_1
XFILLER_98_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09875_ sha256cu.msg_scheduler.mreg_12\[22\] _04153_ _04162_ _04157_ VGND VGND VPWR
+ VPWR _00437_ sky130_fd_sc_hd__o211a_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ sha256cu.m_out_digest.h_in\[6\] sha256cu.m_out_digest.d_in\[6\] VGND VGND
+ VPWR VPWR _03322_ sky130_fd_sc_hd__nor2_1
XFILLER_97_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _03232_ _03234_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__nand2_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_306 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _02323_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__nand2_1
XANTENNA_317 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _02112_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__buf_4
XANTENNA_328 _01558_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_339 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07639_ sha256cu.m_out_digest.b_in\[7\] sha256cu.m_out_digest.a_in\[7\] VGND VGND
+ VPWR VPWR _02262_ sky130_fd_sc_hd__or2_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10650_ _04580_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__buf_2
XFILLER_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09309_ _03786_ _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__nand2_1
X_10581_ sha256cu.msg_scheduler.mreg_9\[28\] _04561_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__or2_1
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12320_ sha256cu.msg_scheduler.mreg_0\[31\] _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ _06028_ _06053_ _06055_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__o21a_1
XFILLER_79_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11202_ sha256cu.m_pad_pars.block_512\[30\]\[4\] _05009_ _04977_ sha256cu.m_pad_pars.block_512\[46\]\[4\]
+ _05056_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__a221o_1
XFILLER_5_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12182_ sha256cu.msg_scheduler.mreg_9\[25\] sha256cu.msg_scheduler.mreg_0\[25\] VGND
+ VGND VPWR VPWR _05990_ sky130_fd_sc_hd__nand2_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11133_ _01940_ _04953_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__or2_1
XFILLER_110_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11064_ _04748_ _01953_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__nor2_1
X_10015_ sha256cu.msg_scheduler.mreg_1\[9\] _04234_ _04244_ _04237_ VGND VGND VPWR
+ VPWR _00501_ sky130_fd_sc_hd__o211a_1
XFILLER_1_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14823_ clknet_leaf_13_clk _01337_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[50\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11966_ _05781_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__or2_1
X_14754_ clknet_leaf_103_clk _01268_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13705_ clknet_leaf_83_clk _00251_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[28\]
+ sky130_fd_sc_hd__dfxtp_4
X_10917_ _04755_ _04766_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__nand2_1
X_14685_ clknet_leaf_122_clk _01199_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11897_ _05688_ _05692_ _05689_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__a21boi_1
X_13636_ clknet_leaf_86_clk _00182_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10848_ _01975_ _04722_ _04723_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__and3_1
X_10779_ sha256cu.msg_scheduler.mreg_11\[17\] _04672_ _04680_ _04675_ VGND VGND VPWR
+ VPWR _00829_ sky130_fd_sc_hd__o211a_1
XFILLER_81_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13567_ clknet_leaf_69_clk _00113_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12518_ _01965_ _04962_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__nand2_2
X_13498_ sha256cu.counter_iteration\[6\] _00053_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__and2b_1
XFILLER_145_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12449_ _06195_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14119_ clknet_leaf_32_clk _00665_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07990_ _02600_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06941_ _01571_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_4
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09660_ sha256cu.m_out_digest.h_in\[24\] _02369_ _02478_ sha256cu.m_out_digest.g_in\[24\]
+ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__o22a_1
XFILLER_95_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08611_ sha256cu.m_out_digest.b_in\[29\] _03177_ _03176_ _02272_ VGND VGND VPWR VPWR
+ _00156_ sky130_fd_sc_hd__o22a_1
X_06872_ sha256cu.msg_scheduler.counter_iteration\[6\] _01566_ VGND VGND VPWR VPWR
+ _01567_ sky130_fd_sc_hd__and2_1
XFILLER_94_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09591_ _02112_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__buf_4
X_08542_ _03101_ _03112_ _03141_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__o21bai_1
XFILLER_63_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08473_ _03037_ _03066_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__or2_1
XFILLER_23_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07424_ sha256cu.m_out_digest.a_in\[14\] sha256cu.m_out_digest.a_in\[3\] VGND VGND
+ VPWR VPWR _02053_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07355_ sha256cu.m_pad_pars.add_out0\[4\] _01976_ _01992_ VGND VGND VPWR VPWR _01993_
+ sky130_fd_sc_hd__and3_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07286_ _01932_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09025_ sha256cu.iter_processing.w\[13\] _02488_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__and2_1
XFILLER_144_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09927_ sha256cu.msg_scheduler.mreg_0\[3\] _04167_ _04194_ _04171_ VGND VGND VPWR
+ VPWR _00463_ sky130_fd_sc_hd__o211a_1
XFILLER_120_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09858_ sha256cu.msg_scheduler.mreg_12\[15\] _04140_ _04152_ _04144_ VGND VGND VPWR
+ VPWR _00430_ sky130_fd_sc_hd__o211a_1
XFILLER_46_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _03304_ _03305_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__xnor2_1
X_09789_ sha256cu.msg_scheduler.mreg_14\[18\] _04106_ VGND VGND VPWR VPWR _04113_
+ sky130_fd_sc_hd__or2_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_125 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ sha256cu.msg_scheduler.mreg_9\[10\] sha256cu.msg_scheduler.mreg_0\[10\] VGND
+ VGND VPWR VPWR _05643_ sky130_fd_sc_hd__nand2_1
XFILLER_61_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_103 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_147 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _05575_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__nor2_1
XANTENNA_158 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_136 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10702_ sha256cu.msg_scheduler.mreg_11\[16\] _04627_ VGND VGND VPWR VPWR _04637_
+ sky130_fd_sc_hd__or2_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_169 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11682_ sha256cu.msg_scheduler.mreg_1\[11\] sha256cu.msg_scheduler.mreg_1\[7\] VGND
+ VGND VPWR VPWR _05511_ sky130_fd_sc_hd__xnor2_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14470_ clknet_leaf_102_clk _00984_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10633_ sha256cu.msg_scheduler.mreg_10\[18\] _04588_ VGND VGND VPWR VPWR _04598_
+ sky130_fd_sc_hd__or2_1
X_13421_ sha256cu.m_pad_pars.block_512\[62\]\[7\] _01928_ VGND VGND VPWR VPWR _06712_
+ sky130_fd_sc_hd__and2_1
XFILLER_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10564_ sha256cu.msg_scheduler.mreg_8\[20\] _04554_ _04558_ _04557_ VGND VGND VPWR
+ VPWR _00736_ sky130_fd_sc_hd__o211a_1
X_13352_ _06676_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12303_ _06103_ _06104_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__or2_1
X_10495_ sha256cu.msg_scheduler.mreg_7\[23\] _04513_ _04518_ _04516_ VGND VGND VPWR
+ VPWR _00707_ sky130_fd_sc_hd__o211a_1
XFILLER_127_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13283_ _06640_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12234_ _06038_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__nor2_1
XFILLER_123_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xpassword_cracker_290 VGND VGND VPWR VPWR password_cracker_290/HI password_count[30]
+ sky130_fd_sc_hd__conb_1
X_12165_ _05941_ _05945_ _05942_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__a21boi_1
XFILLER_107_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11116_ _04973_ _04974_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__nor2_2
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12096_ _05874_ _05879_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__and3_1
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11047_ _04747_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__clkbuf_4
Xinput9 hash[107] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14806_ clknet_leaf_114_clk _01320_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12998_ _06488_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__clkbuf_1
X_11949_ _05764_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_71_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_44_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14737_ clknet_leaf_0_clk _01251_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14668_ clknet_leaf_14_clk _01182_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13619_ clknet_leaf_59_clk _00165_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14599_ clknet_leaf_15_clk _01113_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_07140_ _01644_ _01610_ _01660_ _01797_ _01570_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__a311o_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07071_ _01595_ _01751_ _01596_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__o21a_1
XFILLER_126_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07973_ _02553_ _02554_ _02586_ _02017_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__o31a_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09712_ sha256cu.msg_scheduler.mreg_14\[16\] _04060_ _04069_ _04064_ VGND VGND VPWR
+ VPWR _00367_ sky130_fd_sc_hd__o211a_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06924_ _01611_ _01614_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__or2_2
XFILLER_83_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06855_ _01549_ _01550_ _01551_ _01552_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__or4_1
X_09643_ _02112_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09574_ _02923_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__clkbuf_4
X_08525_ sha256cu.m_out_digest.b_in\[30\] _02304_ _03124_ VGND VGND VPWR VPWR _03125_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06786_ net199 net203 net202 net205 VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__or4_2
XFILLER_36_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08456_ _03040_ _03011_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07407_ _02016_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__buf_4
XFILLER_23_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08387_ _02953_ _02954_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__nand2_1
XFILLER_149_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07338_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07269_ _01911_ _01921_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__or2_1
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10280_ _01972_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__buf_2
X_09008_ _03496_ _03497_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__nand2_1
XFILLER_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13970_ clknet_leaf_54_clk _00516_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[24\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12921_ sha256cu.m_pad_pars.block_512\[33\]\[3\] _06444_ VGND VGND VPWR VPWR _06448_
+ sky130_fd_sc_hd__and2_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ sha256cu.m_pad_pars.block_512\[29\]\[3\] _06407_ VGND VGND VPWR VPWR _06411_
+ sky130_fd_sc_hd__and2_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _05598_ _05602_ _05599_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__a21boi_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _06374_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__clkbuf_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _05557_ _05559_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__or2_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14522_ clknet_leaf_126_clk _01036_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11665_ sha256cu.msg_scheduler.mreg_14\[20\] sha256cu.msg_scheduler.mreg_14\[13\]
+ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__xnor2_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14453_ clknet_leaf_4_clk _00967_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10616_ _04547_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_13404_ _06703_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14384_ clknet_leaf_47_clk _00898_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_11596_ _04698_ _04705_ _02068_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10547_ sha256cu.msg_scheduler.mreg_9\[13\] _04548_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__or2_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13335_ _06667_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__clkbuf_1
X_10478_ sha256cu.msg_scheduler.mreg_8\[16\] _04507_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__or2_1
XFILLER_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13266_ _06631_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
X_12217_ _05996_ _06000_ _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__a21oi_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13197_ sha256cu.m_pad_pars.block_512\[49\]\[4\] _06590_ VGND VGND VPWR VPWR _06595_
+ sky130_fd_sc_hd__and2_1
XFILLER_111_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12148_ _05956_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12079_ _05885_ _05890_ _05891_ _05442_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__o211a_1
XFILLER_84_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_64_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09290_ _03764_ _03768_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__and2_1
X_08310_ _02914_ _02915_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__nand2_1
X_08241_ sha256cu.m_out_digest.a_in\[25\] _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__xnor2_1
XANTENNA_14 _01554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_25 sha256cu.msg_scheduler.mreg_14\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08172_ _02745_ _02779_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__o21ai_1
XANTENNA_58 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07123_ _01584_ _01797_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__or2_1
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07054_ _01636_ _01689_ _00456_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07956_ sha256cu.m_out_digest.h_in\[14\] _02528_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__nand2_1
XFILLER_87_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06907_ sha256cu.iter_processing.rst _01579_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__nand2_4
X_07887_ _02501_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09626_ sha256cu.m_out_digest.g_in\[26\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[26\]
+ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__o22a_1
XFILLER_56_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06838_ net126 net129 net128 net131 VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__or4_1
X_09557_ sha256cu.m_out_digest.f_in\[1\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[1\]
+ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_35_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
X_09488_ _03082_ _03960_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__xor2_1
XFILLER_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08508_ _03068_ _03071_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__nand3_1
XFILLER_24_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08439_ _02198_ sha256cu.m_out_digest.a_in\[9\] VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11450_ sha256cu.m_pad_pars.add_out0\[3\] sha256cu.m_pad_pars.add_out0\[2\] VGND
+ VGND VPWR VPWR _05293_ sky130_fd_sc_hd__and2b_2
X_10401_ sha256cu.msg_scheduler.mreg_6\[14\] _04461_ _04465_ _04464_ VGND VGND VPWR
+ VPWR _00666_ sky130_fd_sc_hd__o211a_1
X_11381_ sha256cu.m_pad_pars.block_512\[5\]\[6\] _05160_ _05165_ sha256cu.m_pad_pars.block_512\[37\]\[6\]
+ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__a221o_1
X_10332_ sha256cu.msg_scheduler.mreg_6\[17\] _04415_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__or2_1
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13120_ sha256cu.m_pad_pars.block_512\[45\]\[0\] _06553_ VGND VGND VPWR VPWR _06554_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13051_ sha256cu.m_pad_pars.block_512\[41\]\[0\] _06516_ VGND VGND VPWR VPWR _06517_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10263_ sha256cu.msg_scheduler.mreg_5\[20\] _04374_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__or2_1
XFILLER_105_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12002_ sha256cu.iter_processing.w\[17\] _05666_ _05817_ _05640_ VGND VGND VPWR VPWR
+ _00915_ sky130_fd_sc_hd__o211a_1
X_10194_ sha256cu.msg_scheduler.mreg_4\[22\] _04335_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__or2_1
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13953_ clknet_leaf_52_clk _00499_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_13884_ clknet_leaf_24_clk _00430_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12904_ _06438_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__clkbuf_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12835_ sha256cu.m_pad_pars.block_512\[28\]\[3\] _06398_ VGND VGND VPWR VPWR _06402_
+ sky130_fd_sc_hd__and2_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14505_ clknet_leaf_16_clk _01019_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _06365_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11717_ _05543_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__or2b_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _06328_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_1
Xinput12 hash[10] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_11648_ _05466_ _05467_ _05478_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__a21o_1
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14436_ clknet_leaf_97_clk _00950_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput23 hash[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput45 hash[13] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
X_14367_ clknet_leaf_77_clk _00881_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput34 hash[12] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
X_11579_ _05414_ _05307_ _04761_ _01952_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__o2bb2a_1
Xinput56 hash[14] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput89 hash[17] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput78 hash[16] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
Xinput67 hash[15] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
X_13318_ _06658_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14298_ clknet_leaf_90_clk _00000_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13249_ _06622_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07810_ _02426_ _02428_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__xnor2_2
XFILLER_111_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08790_ _01972_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__buf_4
X_07741_ _02334_ _02361_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__nand2_1
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07672_ sha256cu.m_out_digest.b_in\[8\] sha256cu.m_out_digest.a_in\[8\] VGND VGND
+ VPWR VPWR _02294_ sky130_fd_sc_hd__or2_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09411_ _03885_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__xor2_1
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_53_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09342_ _03818_ _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__nand2_1
XFILLER_41_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09273_ _03751_ _03753_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__xor2_1
X_08224_ _02829_ _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08155_ _02702_ _02727_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__nor2_1
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07106_ _01743_ _01647_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__nor2_1
X_08086_ _02630_ _02696_ _02697_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__a21oi_2
X_07037_ _01640_ _01719_ _01703_ _01690_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__a22o_1
XFILLER_114_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08988_ _03476_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__nor2_1
X_07939_ _02545_ _02549_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__and2b_1
XFILLER_84_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10950_ _04759_ _04791_ _04816_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__o21bai_2
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09609_ sha256cu.m_out_digest.g_in\[13\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[13\]
+ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__a22o_1
XFILLER_113_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10881_ sha256cu.m_pad_pars.add_512_block\[1\] _01939_ VGND VGND VPWR VPWR _04748_
+ sky130_fd_sc_hd__nand2_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12620_ _06287_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12551_ sha256cu.m_pad_pars.block_512\[11\]\[7\] _04946_ _06249_ VGND VGND VPWR VPWR
+ _06250_ sky130_fd_sc_hd__mux2_1
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11502_ sha256cu.m_pad_pars.block_512\[52\]\[2\] _05310_ _05288_ sha256cu.m_pad_pars.block_512\[48\]\[2\]
+ _05342_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__a221o_1
X_12482_ sha256cu.m_pad_pars.block_512\[7\]\[7\] _04923_ _01983_ VGND VGND VPWR VPWR
+ _06213_ sky130_fd_sc_hd__mux2_1
XFILLER_138_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14221_ clknet_leaf_30_clk _00767_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11433_ _04924_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__nor2_1
XFILLER_153_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14152_ clknet_leaf_32_clk _00698_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11364_ sha256cu.data_in_padd\[20\] _04741_ _04742_ _05210_ VGND VGND VPWR VPWR _00883_
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10315_ sha256cu.msg_scheduler.mreg_5\[9\] _04407_ _04416_ _04410_ VGND VGND VPWR
+ VPWR _00629_ sky130_fd_sc_hd__o211a_1
X_14083_ clknet_leaf_37_clk _00629_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13103_ sha256cu.m_pad_pars.block_512\[44\]\[0\] _06544_ VGND VGND VPWR VPWR _06545_
+ sky130_fd_sc_hd__and2_1
X_11295_ _04819_ _05136_ _05145_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__o21ba_1
X_10246_ sha256cu.msg_scheduler.mreg_4\[12\] _04367_ _04376_ _04370_ VGND VGND VPWR
+ VPWR _00600_ sky130_fd_sc_hd__o211a_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13034_ sha256cu.m_pad_pars.block_512\[40\]\[0\] _06507_ VGND VGND VPWR VPWR _06508_
+ sky130_fd_sc_hd__and2_1
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10177_ sha256cu.msg_scheduler.mreg_3\[14\] _04328_ _04337_ _04331_ VGND VGND VPWR
+ VPWR _00570_ sky130_fd_sc_hd__o211a_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13936_ clknet_leaf_53_clk _00482_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13867_ clknet_leaf_21_clk _00413_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13798_ clknet_leaf_81_clk _00344_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12818_ sha256cu.m_pad_pars.block_512\[27\]\[3\] _06389_ VGND VGND VPWR VPWR _06393_
+ sky130_fd_sc_hd__and2_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _06356_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14419_ clknet_leaf_107_clk _00933_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_512_block\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09960_ sha256cu.msg_scheduler.mreg_0\[17\] _04208_ _04213_ _04211_ VGND VGND VPWR
+ VPWR _00477_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_6_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
X_08911_ sha256cu.iter_processing.w\[9\] _02338_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__or2_1
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09891_ sha256cu.msg_scheduler.mreg_13\[29\] _04160_ VGND VGND VPWR VPWR _04172_
+ sky130_fd_sc_hd__or2_1
XFILLER_58_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__nand2_1
XFILLER_112_774 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ sha256cu.K\[4\] VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__inv_2
XFILLER_97_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07724_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__inv_2
X_07655_ sha256cu.m_out_digest.h_in\[6\] _02235_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__nand2_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07586_ _02172_ _02170_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__and2b_1
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ _03802_ _03803_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__nor2_1
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09256_ sha256cu.iter_processing.w\[21\] _02785_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__nor2_1
X_08207_ _02775_ _02813_ _02814_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__o21a_1
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09187_ _03647_ _03648_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__nor2_1
XFILLER_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08138_ _02745_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08069_ sha256cu.m_out_digest.h_in\[17\] _02646_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__nand2_1
XFILLER_150_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10100_ sha256cu.msg_scheduler.mreg_2\[13\] _04288_ _04293_ _04291_ VGND VGND VPWR
+ VPWR _00537_ sky130_fd_sc_hd__o211a_1
XFILLER_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11080_ _04799_ _04936_ _04939_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__a21bo_1
XFILLER_1_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10031_ sha256cu.msg_scheduler.mreg_1\[16\] _04247_ _04253_ _04250_ VGND VGND VPWR
+ VPWR _00508_ sky130_fd_sc_hd__o211a_1
Xinput202 hash[50] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput224 hash[70] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
Xinput235 hash[80] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__buf_2
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput213 hash[60] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput257 reset VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput246 hash[90] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14770_ clknet_leaf_2_clk _01284_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13721_ clknet_leaf_65_clk _00267_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11982_ sha256cu.msg_scheduler.mreg_9\[17\] sha256cu.msg_scheduler.mreg_0\[17\] VGND
+ VGND VPWR VPWR _05798_ sky130_fd_sc_hd__or2_1
XFILLER_72_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10933_ _04795_ _04797_ _04799_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__and3b_2
XFILLER_44_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13652_ clknet_4_15_0_clk _00198_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10864_ sha256cu.m_pad_pars.add_out3\[5\] VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__inv_2
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ clknet_leaf_73_clk _00129_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10795_ sha256cu.msg_scheduler.mreg_11\[24\] _04685_ _04689_ _04688_ VGND VGND VPWR
+ VPWR _00836_ sky130_fd_sc_hd__o211a_1
X_12603_ _06278_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _02068_ sha256cu.m_pad_pars.block_512\[10\]\[7\] _06240_ VGND VGND VPWR VPWR
+ _01024_ sky130_fd_sc_hd__a21o_1
XFILLER_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12465_ sha256cu.m_pad_pars.block_512\[6\]\[7\] _05099_ _01983_ VGND VGND VPWR VPWR
+ _06204_ sky130_fd_sc_hd__mux2_1
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14204_ clknet_leaf_45_clk _00750_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12396_ _06167_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__clkbuf_1
X_11416_ _04769_ _05129_ _05259_ sha256cu.m_pad_pars.block_512\[9\]\[7\] VGND VGND
+ VPWR VPWR _05260_ sky130_fd_sc_hd__o22a_1
X_14135_ clknet_leaf_34_clk _00681_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11347_ sha256cu.m_pad_pars.block_512\[61\]\[3\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[3\]
+ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__a22o_1
XFILLER_125_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14066_ clknet_leaf_38_clk _00612_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11278_ _01941_ _04749_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__or2_2
X_10229_ sha256cu.msg_scheduler.mreg_4\[5\] _04354_ _04366_ _04357_ VGND VGND VPWR
+ VPWR _00593_ sky130_fd_sc_hd__o211a_1
X_13017_ sha256cu.m_pad_pars.block_512\[39\]\[0\] _06498_ VGND VGND VPWR VPWR _06499_
+ sky130_fd_sc_hd__and2_1
XFILLER_121_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13919_ clknet_leaf_44_clk _00465_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14899_ clknet_leaf_1_clk _01413_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_07440_ sha256cu.m_out_digest.a_in\[1\] _02040_ _02067_ _02068_ VGND VGND VPWR VPWR
+ _00096_ sky130_fd_sc_hd__a211o_1
XFILLER_50_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07371_ sha256cu.counter_iteration\[0\] _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__nand2_1
XFILLER_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09110_ sha256cu.K\[16\] _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09041_ sha256cu.m_out_digest.e_in\[13\] _02440_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__or2_1
XFILLER_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09943_ sha256cu.msg_scheduler.mreg_1\[10\] _04202_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__or2_1
XFILLER_100_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09874_ sha256cu.msg_scheduler.mreg_13\[22\] _04160_ VGND VGND VPWR VPWR _04162_
+ sky130_fd_sc_hd__or2_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ sha256cu.K\[6\] _03320_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _03240_ _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_307 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _02324_ _02325_ _02326_ _02328_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__a211oi_4
XANTENNA_318 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08687_ sha256cu.m_out_digest.d_in\[29\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[29\]
+ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__o22a_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07638_ sha256cu.iter_processing.w\[6\] _02226_ _02225_ VGND VGND VPWR VPWR _02261_
+ sky130_fd_sc_hd__a21o_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07569_ sha256cu.iter_processing.w\[5\] _02193_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09308_ sha256cu.m_out_digest.h_in\[23\] sha256cu.m_out_digest.d_in\[23\] VGND VGND
+ VPWR VPWR _03787_ sky130_fd_sc_hd__nand2_1
XFILLER_22_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10580_ _04447_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__buf_2
X_09239_ _03664_ _03691_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__nand2_1
XFILLER_6_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12250_ _06024_ _06045_ _06047_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12181_ sha256cu.msg_scheduler.mreg_9\[25\] sha256cu.msg_scheduler.mreg_0\[25\] VGND
+ VGND VPWR VPWR _05989_ sky130_fd_sc_hd__or2_1
XFILLER_108_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11201_ sha256cu.m_pad_pars.block_512\[10\]\[4\] _04963_ _05051_ _05055_ VGND VGND
+ VPWR VPWR _05056_ sky130_fd_sc_hd__a211o_1
X_11132_ _04990_ _04967_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__nand2_2
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11063_ sha256cu.m_pad_pars.block_512\[7\]\[7\] _04922_ _04772_ VGND VGND VPWR VPWR
+ _04923_ sky130_fd_sc_hd__o21a_1
X_10014_ sha256cu.msg_scheduler.mreg_2\[9\] _04241_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__or2_1
XFILLER_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14822_ clknet_leaf_102_clk _01336_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11965_ _05755_ _05759_ _05756_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__a21boi_2
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14753_ clknet_leaf_106_clk _01267_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13704_ clknet_leaf_83_clk _00250_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[27\]
+ sky130_fd_sc_hd__dfxtp_4
X_10916_ sha256cu.m_pad_pars.block_512\[27\]\[0\] _04757_ _04765_ sha256cu.m_pad_pars.block_512\[3\]\[0\]
+ _04782_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__a221o_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14684_ clknet_leaf_122_clk _01198_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11896_ _05713_ _05715_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__xor2_1
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13635_ clknet_leaf_87_clk _00181_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10847_ _01980_ _04720_ _04721_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__or3b_1
XFILLER_20_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10778_ sha256cu.msg_scheduler.mreg_12\[17\] _04679_ VGND VGND VPWR VPWR _04680_
+ sky130_fd_sc_hd__or2_1
X_13566_ clknet_leaf_69_clk _00112_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12517_ _06231_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13497_ _06762_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12448_ sha256cu.m_pad_pars.block_512\[5\]\[7\] _05238_ _01983_ VGND VGND VPWR VPWR
+ _06195_ sky130_fd_sc_hd__mux2_1
XFILLER_5_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12379_ sha256cu.m_pad_pars.block_512\[1\]\[6\] _06152_ VGND VGND VPWR VPWR _06159_
+ sky130_fd_sc_hd__and2_1
X_14118_ clknet_leaf_32_clk _00664_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14049_ clknet_leaf_40_clk _00595_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_06940_ _00457_ _01599_ _01619_ _01630_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__a2bb2o_1
X_06871_ sha256cu.msg_scheduler.counter_iteration\[5\] sha256cu.msg_scheduler.counter_iteration\[4\]
+ _01565_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__nor3_4
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08610_ sha256cu.m_out_digest.b_in\[28\] _03177_ _03176_ _02232_ VGND VGND VPWR VPWR
+ _00155_ sky130_fd_sc_hd__o22a_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09590_ sha256cu.m_out_digest.f_in\[29\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[29\]
+ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__a22o_1
X_08541_ sha256cu.K\[30\] _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__xor2_1
X_08472_ _02232_ _03031_ _03071_ _03073_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__a22o_1
X_07423_ _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__inv_2
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07354_ sha256cu.m_pad_pars.add_out0\[3\] sha256cu.m_pad_pars.add_out0\[2\] VGND
+ VGND VPWR VPWR _01992_ sky130_fd_sc_hd__and2_2
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07285_ sha256cu.m_pad_pars.m_size\[6\] sha256cu.m_pad_pars.block_512\[63\]\[6\]
+ _01923_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__mux2_1
X_09024_ sha256cu.iter_processing.w\[13\] _02488_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__nor2_1
XFILLER_144_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09926_ sha256cu.msg_scheduler.mreg_1\[3\] _04174_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__or2_1
XFILLER_98_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09857_ sha256cu.msg_scheduler.mreg_13\[15\] _04147_ VGND VGND VPWR VPWR _04152_
+ sky130_fd_sc_hd__or2_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08808_ _03271_ _03274_ _03273_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__o21ai_1
X_09788_ _04044_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__buf_2
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _03237_ _03238_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__nor2_1
XFILLER_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_104 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_148 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11750_ _05550_ _05554_ _05551_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__a21boi_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10701_ sha256cu.msg_scheduler.mreg_10\[15\] _04633_ _04635_ _04636_ VGND VGND VPWR
+ VPWR _00795_ sky130_fd_sc_hd__o211a_1
XANTENNA_159 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _05508_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__nand2_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10632_ sha256cu.msg_scheduler.mreg_9\[17\] _04594_ _04596_ _04597_ VGND VGND VPWR
+ VPWR _00765_ sky130_fd_sc_hd__o211a_1
X_13420_ _06711_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__clkbuf_1
X_10563_ sha256cu.msg_scheduler.mreg_9\[20\] _04548_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__or2_1
X_13351_ sha256cu.m_pad_pars.block_512\[58\]\[5\] _06671_ VGND VGND VPWR VPWR _06676_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12302_ _06103_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nand2_1
XFILLER_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10494_ sha256cu.msg_scheduler.mreg_8\[23\] _04507_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__or2_1
X_13282_ sha256cu.m_pad_pars.block_512\[54\]\[4\] _06635_ VGND VGND VPWR VPWR _06640_
+ sky130_fd_sc_hd__and2_1
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12233_ _06010_ _06014_ _06011_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__a21boi_1
Xpassword_cracker_280 VGND VGND VPWR VPWR password_cracker_280/HI password_count[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12164_ _05970_ _05972_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__xor2_1
Xpassword_cracker_291 VGND VGND VPWR VPWR password_cracker_291/HI password_count[31]
+ sky130_fd_sc_hd__conb_1
X_12095_ _05904_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11115_ _04701_ _04779_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__nor2_1
X_11046_ sha256cu.m_pad_pars.block_512\[55\]\[7\] _04833_ _04905_ _04738_ VGND VGND
+ VPWR VPWR _04906_ sky130_fd_sc_hd__a22o_1
XFILLER_49_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14805_ clknet_leaf_4_clk _01319_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12997_ sha256cu.m_pad_pars.block_512\[37\]\[7\] _05247_ _06442_ VGND VGND VPWR VPWR
+ _06488_ sky130_fd_sc_hd__mux2_1
X_14736_ clknet_leaf_4_clk _01250_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11948_ sha256cu.msg_scheduler.mreg_14\[25\] _05765_ VGND VGND VPWR VPWR _05766_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_44_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11879_ _05697_ _05699_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__nand2_1
X_14667_ clknet_leaf_13_clk _01181_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13618_ clknet_leaf_59_clk _00164_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14598_ clknet_leaf_102_clk _01112_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13549_ clknet_leaf_74_clk _00095_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_71_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07070_ _01606_ _01750_ _01639_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__a21oi_2
XFILLER_146_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07972_ _02553_ _02554_ _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__o21ai_1
X_09711_ sha256cu.iter_processing.w\[16\] _04067_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__or2_1
XFILLER_19_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06923_ _01586_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__or2_1
X_09642_ sha256cu.m_out_digest.h_in\[8\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[8\]
+ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__o22a_1
X_06854_ net37 net40 net39 net42 VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__or4_4
XFILLER_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09573_ sha256cu.m_out_digest.f_in\[14\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[14\]
+ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__o22a_1
XFILLER_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06785_ net191 net194 net193 net196 VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__or4_4
X_08524_ sha256cu.m_out_digest.b_in\[30\] _02304_ sha256cu.m_out_digest.c_in\[30\]
+ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__a21o_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08455_ _03055_ _03056_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__nand2_1
XFILLER_23_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07406_ sha256cu.K\[0\] _02034_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__or2_1
X_08386_ _02953_ _02954_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__nor2_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07337_ _01911_ _01961_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__nor2_1
XFILLER_51_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07268_ _01920_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__clkbuf_4
X_09007_ _03493_ _03495_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__or2_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07199_ _01644_ _01862_ _01863_ _01571_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__o211a_1
XFILLER_144_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09909_ sha256cu.msg_scheduler.counter_iteration\[4\] _04181_ VGND VGND VPWR VPWR
+ _04184_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12920_ _06447_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12851_ _06410_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11802_ _05623_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__xor2_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ sha256cu.m_pad_pars.block_512\[25\]\[2\] _06371_ VGND VGND VPWR VPWR _06374_
+ sky130_fd_sc_hd__and2_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _05557_ _05559_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nand2_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14521_ clknet_leaf_126_clk _01035_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11664_ _05492_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__and2_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ clknet_leaf_5_clk _00966_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10615_ sha256cu.msg_scheduler.mreg_9\[10\] _04581_ _04587_ _04584_ VGND VGND VPWR
+ VPWR _00758_ sky130_fd_sc_hd__o211a_1
X_13403_ sha256cu.m_pad_pars.block_512\[61\]\[6\] _06693_ VGND VGND VPWR VPWR _06703_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11595_ _05429_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
X_14383_ clknet_leaf_107_clk _00897_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.temp_chk
+ sky130_fd_sc_hd__dfxtp_1
X_10546_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__clkbuf_2
XFILLER_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13334_ sha256cu.m_pad_pars.block_512\[57\]\[5\] _06660_ VGND VGND VPWR VPWR _06667_
+ sky130_fd_sc_hd__and2_1
X_10477_ sha256cu.msg_scheduler.mreg_7\[15\] _04500_ _04508_ _04503_ VGND VGND VPWR
+ VPWR _00699_ sky130_fd_sc_hd__o211a_1
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13265_ sha256cu.m_pad_pars.block_512\[53\]\[4\] _06626_ VGND VGND VPWR VPWR _06631_
+ sky130_fd_sc_hd__and2_1
XFILLER_108_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12216_ _06021_ _06022_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__nand2_1
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13196_ _06594_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12147_ _05934_ _05937_ _05931_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12078_ _05885_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__nand2_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11029_ sha256cu.m_pad_pars.block_512\[15\]\[5\] _04781_ _04800_ sha256cu.m_pad_pars.block_512\[39\]\[5\]
+ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__a22o_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14719_ clknet_leaf_100_clk _01233_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[37\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08240_ _02027_ sha256cu.m_out_digest.a_in\[4\] VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__xnor2_2
XANTENNA_26 sha256cu.msg_scheduler.mreg_9\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ sha256cu.m_out_digest.h_in\[20\] _02744_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__nand2_1
XANTENNA_15 _01554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07122_ _01719_ _01673_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__nor2_1
XFILLER_146_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07053_ _01648_ _01687_ _01733_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__a31o_1
XFILLER_99_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07955_ _02566_ _02569_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__xnor2_2
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06906_ _01581_ _01585_ _01591_ _01595_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__o32a_1
X_07886_ _02448_ _02458_ _02502_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__o21ba_1
X_09625_ sha256cu.m_out_digest.g_in\[25\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[25\]
+ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__o22a_1
XFILLER_44_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06837_ net121 net125 net124 net127 VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__or4_1
X_09556_ sha256cu.m_out_digest.f_in\[0\] _03559_ _03192_ sha256cu.m_out_digest.e_in\[0\]
+ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__a22o_1
X_09487_ _03958_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__nand2_1
XFILLER_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08507_ _03105_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__nand2_1
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08438_ _03002_ _03004_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__nand2_1
XFILLER_11_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08369_ sha256cu.iter_processing.w\[26\] _02972_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__xor2_1
X_10400_ sha256cu.msg_scheduler.mreg_7\[14\] _04455_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__or2_1
XFILLER_125_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11380_ sha256cu.m_pad_pars.block_512\[53\]\[6\] _05161_ _05224_ _05024_ VGND VGND
+ VPWR VPWR _05225_ sky130_fd_sc_hd__a22o_1
XFILLER_20_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10331_ sha256cu.msg_scheduler.mreg_5\[16\] _04421_ _04425_ _04424_ VGND VGND VPWR
+ VPWR _00636_ sky130_fd_sc_hd__o211a_1
XFILLER_109_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10262_ sha256cu.msg_scheduler.mreg_4\[19\] _04380_ _04385_ _04383_ VGND VGND VPWR
+ VPWR _00607_ sky130_fd_sc_hd__o211a_1
XFILLER_118_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13050_ _01986_ _05131_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__or2_2
XFILLER_140_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12001_ sha256cu.data_in_padd\[17\] _05667_ _05816_ _05445_ VGND VGND VPWR VPWR _05817_
+ sky130_fd_sc_hd__a211o_1
X_10193_ sha256cu.msg_scheduler.mreg_3\[21\] _04341_ _04346_ _04344_ VGND VGND VPWR
+ VPWR _00577_ sky130_fd_sc_hd__o211a_1
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13952_ clknet_leaf_54_clk _00498_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12903_ sha256cu.m_pad_pars.block_512\[32\]\[3\] _06434_ VGND VGND VPWR VPWR _06438_
+ sky130_fd_sc_hd__and2_1
XFILLER_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13883_ clknet_leaf_24_clk _00429_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12834_ _06401_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12765_ sha256cu.m_pad_pars.block_512\[24\]\[2\] _06362_ VGND VGND VPWR VPWR _06365_
+ sky130_fd_sc_hd__and2_1
XFILLER_15_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _05515_ _05529_ _05542_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__a21o_1
X_14504_ clknet_leaf_8_clk _01018_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ sha256cu.m_pad_pars.block_512\[20\]\[2\] _06325_ VGND VGND VPWR VPWR _06328_
+ sky130_fd_sc_hd__and2_1
X_11647_ _05475_ _05477_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__xnor2_1
Xinput13 hash[110] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlymetal6s2s_1
X_14435_ clknet_leaf_96_clk _00949_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput46 hash[140] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
X_14366_ clknet_leaf_77_clk _00880_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput35 hash[130] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 hash[120] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
X_11578_ sha256cu.m_pad_pars.block_512\[52\]\[7\] VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__inv_1
Xinput57 hash[150] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
X_10529_ sha256cu.msg_scheduler.mreg_9\[6\] _04534_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__or2_1
XFILLER_116_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput68 hash[160] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
X_13317_ sha256cu.m_pad_pars.block_512\[56\]\[5\] _01924_ VGND VGND VPWR VPWR _06658_
+ sky130_fd_sc_hd__and2_1
Xinput79 hash[170] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
XFILLER_115_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14297_ clknet_leaf_20_clk _00843_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_13248_ sha256cu.m_pad_pars.block_512\[52\]\[4\] _06617_ VGND VGND VPWR VPWR _06622_
+ sky130_fd_sc_hd__and2_1
X_13179_ sha256cu.m_pad_pars.block_512\[48\]\[4\] _06580_ VGND VGND VPWR VPWR _06585_
+ sky130_fd_sc_hd__and2_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07740_ sha256cu.K\[9\] _02360_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07671_ sha256cu.iter_processing.w\[7\] _02266_ _02265_ VGND VGND VPWR VPWR _02293_
+ sky130_fd_sc_hd__a21o_1
XFILLER_65_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09410_ sha256cu.K\[25\] _03851_ _03853_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__a21o_1
XFILLER_80_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09341_ _03816_ _03817_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__nand2_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09272_ _03719_ _03752_ _03717_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__a21bo_1
XFILLER_60_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08223_ sha256cu.iter_processing.w\[21\] _02786_ _02830_ VGND VGND VPWR VPWR _02831_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_21_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08154_ _02702_ _02727_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__nand2_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08085_ _02619_ _02660_ _02659_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__o21ba_1
X_07105_ _01644_ _01688_ _01779_ _01780_ _01781_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__o32a_1
X_07036_ _01578_ _01625_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__nand2_2
XFILLER_122_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08987_ sha256cu.m_out_digest.h_in\[12\] sha256cu.m_out_digest.d_in\[12\] VGND VGND
+ VPWR VPWR _03477_ sky130_fd_sc_hd__and2_1
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07938_ _02542_ _02544_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__and2b_1
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07869_ sha256cu.m_out_digest.b_in\[13\] _02027_ sha256cu.m_out_digest.c_in\[13\]
+ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__a21o_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09608_ sha256cu.m_out_digest.g_in\[12\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[12\]
+ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__o22a_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10880_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__buf_4
X_09539_ _04007_ _04009_ _04010_ _02068_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__a211o_1
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12550_ _01964_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__buf_4
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12481_ _06212_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__clkbuf_1
X_11501_ sha256cu.m_pad_pars.block_512\[28\]\[2\] _05296_ _05341_ _01921_ VGND VGND
+ VPWR VPWR _05342_ sky130_fd_sc_hd__a22o_1
X_14220_ clknet_leaf_30_clk _00766_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11432_ _04701_ _05129_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__nor2_2
X_14151_ clknet_leaf_31_clk _00697_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13102_ _02111_ _04917_ _05295_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__or3_2
X_11363_ _05202_ _05204_ _05209_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__or3_1
XFILLER_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10314_ sha256cu.msg_scheduler.mreg_6\[9\] _04415_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__or2_1
X_14082_ clknet_leaf_38_clk _00628_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11294_ _04705_ _04792_ _04993_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__nor3_1
X_10245_ sha256cu.msg_scheduler.mreg_5\[12\] _04374_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__or2_1
XFILLER_105_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _06270_ _05319_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__nand2_2
X_10176_ sha256cu.msg_scheduler.mreg_4\[14\] _04335_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__or2_1
XFILLER_120_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13935_ clknet_leaf_52_clk _00481_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13866_ clknet_leaf_21_clk _00412_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12817_ _06392_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13797_ clknet_leaf_88_clk _00343_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ sha256cu.m_pad_pars.block_512\[23\]\[2\] _06353_ VGND VGND VPWR VPWR _06356_
+ sky130_fd_sc_hd__and2_1
XFILLER_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12679_ sha256cu.m_pad_pars.block_512\[19\]\[2\] _06316_ VGND VGND VPWR VPWR _06319_
+ sky130_fd_sc_hd__and2_1
X_14418_ clknet_leaf_106_clk _00932_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_512_block\[2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14349_ clknet_leaf_110_clk _00863_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08910_ _03401_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__or2b_1
XFILLER_143_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09890_ sha256cu.msg_scheduler.mreg_12\[28\] _04167_ _04170_ _04171_ VGND VGND VPWR
+ VPWR _00443_ sky130_fd_sc_hd__o211a_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _03333_ _03335_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__or2_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _03268_ _03269_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__xnor2_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07723_ sha256cu.m_out_digest.e_in\[20\] _02343_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__xnor2_4
XFILLER_84_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07654_ _02271_ _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07585_ _02187_ _02209_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09324_ _03762_ _03769_ _03801_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__nor3_1
XFILLER_34_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09255_ _03734_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__or2_1
X_08206_ sha256cu.m_out_digest.h_in\[21\] _02774_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__nand2_1
X_09186_ _03659_ _03660_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__nand2_1
X_08137_ sha256cu.m_out_digest.e_in\[31\] _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__xnor2_4
XFILLER_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08068_ _02676_ _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07019_ _01702_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__nand2_1
X_10030_ sha256cu.msg_scheduler.mreg_2\[16\] _04241_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__or2_1
XFILLER_88_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput214 hash[61] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
XFILLER_130_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput236 hash[81] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
Xinput225 hash[71] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput203 hash[51] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_124_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput247 hash[91] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
X_11981_ sha256cu.iter_processing.w\[16\] _05666_ _05797_ _05640_ VGND VGND VPWR VPWR
+ _00914_ sky130_fd_sc_hd__o211a_1
X_13720_ clknet_leaf_65_clk _00266_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10932_ _04767_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__and2_1
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13651_ clknet_leaf_59_clk _00197_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10863_ _04734_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ clknet_leaf_73_clk _00128_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10794_ sha256cu.msg_scheduler.mreg_12\[24\] _04679_ VGND VGND VPWR VPWR _04689_
+ sky130_fd_sc_hd__or2_1
X_12602_ sha256cu.m_pad_pars.block_512\[14\]\[6\] _06271_ VGND VGND VPWR VPWR _06278_
+ sky130_fd_sc_hd__and2_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ sha256cu.m_pad_pars.block_512\[10\]\[7\] _05090_ _05091_ _01975_ VGND VGND
+ VPWR VPWR _06240_ sky130_fd_sc_hd__o211a_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14203_ clknet_leaf_45_clk _00749_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12464_ _06203_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12395_ sha256cu.m_pad_pars.block_512\[2\]\[6\] _06160_ VGND VGND VPWR VPWR _06167_
+ sky130_fd_sc_hd__and2_1
X_11415_ _04702_ _05091_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__nor2_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14134_ clknet_leaf_34_clk _00680_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11346_ sha256cu.m_pad_pars.block_512\[29\]\[3\] _05141_ _05135_ sha256cu.m_pad_pars.block_512\[1\]\[3\]
+ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__a221o_1
XFILLER_153_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14065_ clknet_leaf_39_clk _00611_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13016_ _04795_ _04970_ _01972_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__o21ai_4
X_11277_ _04933_ _05124_ _05127_ _01977_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__o211a_2
X_10228_ sha256cu.msg_scheduler.mreg_5\[5\] _04361_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__or2_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10159_ sha256cu.msg_scheduler.mreg_4\[7\] _04322_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__or2_1
XFILLER_94_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13918_ clknet_leaf_44_clk _00464_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14898_ clknet_leaf_1_clk _01412_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13849_ clknet_leaf_21_clk _00395_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07370_ sha256cu.counter_iteration\[3\] sha256cu.counter_iteration\[2\] sha256cu.counter_iteration\[1\]
+ _02004_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__nor4_4
X_09040_ _03496_ _03503_ _03527_ _02065_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__a31o_1
XFILLER_132_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09942_ sha256cu.msg_scheduler.mreg_0\[9\] _04195_ _04203_ _04198_ VGND VGND VPWR
+ VPWR _00469_ sky130_fd_sc_hd__o211a_1
XFILLER_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09873_ sha256cu.msg_scheduler.mreg_12\[21\] _04153_ _04161_ _04157_ VGND VGND VPWR
+ VPWR _00436_ sky130_fd_sc_hd__o211a_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08824_ _03318_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__nor2_1
XFILLER_100_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _03251_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _02260_ _02289_ _02327_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_319 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ sha256cu.m_out_digest.d_in\[28\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[28\]
+ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__a22o_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07637_ sha256cu.K\[6\] _02248_ _02259_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__a21oi_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07568_ _02191_ _02192_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__and2b_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09307_ sha256cu.m_out_digest.h_in\[23\] sha256cu.m_out_digest.d_in\[23\] VGND VGND
+ VPWR VPWR _03786_ sky130_fd_sc_hd__or2_1
X_07499_ sha256cu.m_out_digest.e_in\[28\] _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__xnor2_2
XFILLER_21_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09238_ _03608_ _03637_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__nand2_1
X_09169_ sha256cu.K\[18\] _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12180_ _05977_ _05978_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__or2b_1
XFILLER_79_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11200_ sha256cu.m_pad_pars.block_512\[6\]\[4\] _04957_ _05053_ _05054_ VGND VGND
+ VPWR VPWR _05055_ sky130_fd_sc_hd__a211o_1
XFILLER_150_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11131_ sha256cu.m_pad_pars.add_out2\[3\] sha256cu.m_pad_pars.add_out2\[2\] VGND
+ VGND VPWR VPWR _04990_ sky130_fd_sc_hd__nor2_2
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11062_ _04770_ _04787_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__nor2_1
X_10013_ sha256cu.msg_scheduler.mreg_1\[8\] _04234_ _04243_ _04237_ VGND VGND VPWR
+ VPWR _00500_ sky130_fd_sc_hd__o211a_1
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14821_ clknet_leaf_98_clk _01335_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ _05778_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__xor2_1
X_14752_ clknet_leaf_106_clk _01266_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11895_ sha256cu.msg_scheduler.mreg_1\[31\] _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__xnor2_1
X_13703_ clknet_leaf_83_clk _00249_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[26\]
+ sky130_fd_sc_hd__dfxtp_4
X_10915_ sha256cu.m_pad_pars.block_512\[7\]\[0\] _04774_ _04781_ sha256cu.m_pad_pars.block_512\[15\]\[0\]
+ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a22o_1
XFILLER_44_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14683_ clknet_leaf_121_clk _01197_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10846_ sha256cu.m_pad_pars.add_out2\[3\] sha256cu.m_pad_pars.add_out2\[2\] _01976_
+ _04721_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__a31o_1
X_13634_ clknet_leaf_86_clk _00180_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10777_ _01566_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__clkbuf_2
X_13565_ clknet_leaf_69_clk _00111_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12516_ sha256cu.m_pad_pars.block_512\[9\]\[7\] _05260_ _01983_ VGND VGND VPWR VPWR
+ _06231_ sky130_fd_sc_hd__mux2_1
XFILLER_9_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13496_ _01975_ _06761_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__and2_1
XFILLER_67_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12447_ _06194_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14117_ clknet_leaf_37_clk _00663_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12378_ _06158_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11329_ sha256cu.m_pad_pars.block_512\[9\]\[1\] _05144_ _05147_ sha256cu.m_pad_pars.block_512\[33\]\[1\]
+ _05178_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__a221o_1
X_14048_ clknet_leaf_39_clk _00594_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06870_ sha256cu.msg_scheduler.counter_iteration\[0\] sha256cu.msg_scheduler.counter_iteration\[3\]
+ sha256cu.msg_scheduler.counter_iteration\[2\] sha256cu.msg_scheduler.counter_iteration\[1\]
+ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__or4_2
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08540_ _03138_ _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__or2b_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08471_ _02478_ _03072_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__nor2_1
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07422_ sha256cu.m_out_digest.e_in\[26\] _02050_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__xnor2_2
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07353_ sha256cu.m_pad_pars.add_out0\[3\] _01989_ _01991_ _01971_ _01974_ VGND VGND
+ VPWR VPWR _00086_ sky130_fd_sc_hd__o221a_1
X_07284_ _01931_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09023_ _03510_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09925_ sha256cu.msg_scheduler.mreg_0\[2\] _04167_ _04193_ _04171_ VGND VGND VPWR
+ VPWR _00462_ sky130_fd_sc_hd__o211a_1
XFILLER_131_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09856_ sha256cu.msg_scheduler.mreg_12\[14\] _04140_ _04151_ _04144_ VGND VGND VPWR
+ VPWR _00429_ sky130_fd_sc_hd__o211a_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _03301_ _03303_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09787_ sha256cu.msg_scheduler.mreg_13\[17\] _04099_ _04111_ _04103_ VGND VGND VPWR
+ VPWR _00400_ sky130_fd_sc_hd__o211a_1
X_06999_ _01607_ _01600_ _01602_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__and3_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _03220_ _03218_ _03236_ _02065_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__a31o_1
XFILLER_54_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_116 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_149 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08669_ sha256cu.m_out_digest.d_in\[13\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[13\]
+ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__o22a_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_138 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10700_ _04529_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__buf_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11680_ sha256cu.msg_scheduler.mreg_9\[4\] sha256cu.msg_scheduler.mreg_0\[4\] VGND
+ VGND VPWR VPWR _05509_ sky130_fd_sc_hd__nand2_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10631_ _04529_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__buf_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10562_ sha256cu.msg_scheduler.mreg_8\[19\] _04554_ _04556_ _04557_ VGND VGND VPWR
+ VPWR _00735_ sky130_fd_sc_hd__o211a_1
X_13350_ _06675_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12301_ sha256cu.msg_scheduler.mreg_14\[17\] sha256cu.msg_scheduler.mreg_14\[15\]
+ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__xor2_1
X_13281_ _06639_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
X_10493_ sha256cu.msg_scheduler.mreg_7\[22\] _04513_ _04517_ _04516_ VGND VGND VPWR
+ VPWR _00706_ sky130_fd_sc_hd__o211a_1
X_12232_ _06035_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__xor2_1
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpassword_cracker_270 VGND VGND VPWR VPWR password_cracker_270/HI password_count[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_107_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpassword_cracker_281 VGND VGND VPWR VPWR password_cracker_281/HI password_count[21]
+ sky130_fd_sc_hd__conb_1
XFILLER_122_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12163_ sha256cu.msg_scheduler.mreg_1\[31\] _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12094_ sha256cu.msg_scheduler.mreg_14\[31\] _05905_ VGND VGND VPWR VPWR _05906_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_1_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11114_ _04776_ _04953_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__nor2_2
XFILLER_104_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11045_ sha256cu.m_pad_pars.m_size\[7\] sha256cu.m_pad_pars.block_512\[63\]\[7\]
+ _01921_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__mux2_1
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12996_ _06487_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__clkbuf_1
X_14804_ clknet_leaf_1_clk _01318_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11947_ sha256cu.msg_scheduler.mreg_14\[2\] sha256cu.msg_scheduler.mreg_14\[0\] VGND
+ VGND VPWR VPWR _05765_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14735_ clknet_leaf_4_clk _01249_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[39\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11878_ sha256cu.msg_scheduler.mreg_14\[31\] _05698_ VGND VGND VPWR VPWR _05699_
+ sky130_fd_sc_hd__xnor2_1
X_14666_ clknet_leaf_12_clk _01180_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13617_ clknet_leaf_51_clk _00163_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14597_ clknet_leaf_98_clk _01111_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10829_ sha256cu.m_pad_pars.m_size\[7\] _04706_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__or2_1
X_13548_ clknet_leaf_80_clk _00094_ VGND VGND VPWR VPWR sha256cu.iter_processing.temp_case
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13479_ sha256cu.K\[18\] _06714_ _06719_ _00045_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__a22o_1
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07971_ _02584_ _02585_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__nor2_1
XFILLER_102_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09710_ sha256cu.msg_scheduler.mreg_14\[15\] _04060_ _04068_ _04064_ VGND VGND VPWR
+ VPWR _00366_ sky130_fd_sc_hd__o211a_1
X_06922_ _01589_ _01612_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__nand2_1
X_09641_ sha256cu.m_out_digest.h_in\[7\] _04037_ _04036_ sha256cu.m_out_digest.g_in\[7\]
+ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__a22o_1
XFILLER_110_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06853_ net32 net36 net35 net38 VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__or4_2
X_09572_ sha256cu.m_out_digest.f_in\[13\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[13\]
+ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__o22a_1
X_06784_ net195 net198 net197 net200 VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__or4_1
X_08523_ _03120_ _03122_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__xor2_1
XFILLER_70_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08454_ _03049_ _03054_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__or2_1
X_07405_ sha256cu.K\[0\] _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nand2_1
X_08385_ _02920_ _02955_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__or2_1
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07336_ _01976_ _01977_ sha256cu.m_pad_pars.add_out1\[4\] VGND VGND VPWR VPWR _01978_
+ sky130_fd_sc_hd__a21o_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09006_ _03493_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__nand2_1
X_07267_ _01919_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__buf_4
XFILLER_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07198_ _01584_ _01849_ _01658_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__or3_1
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09908_ _04183_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09839_ sha256cu.msg_scheduler.mreg_13\[7\] _04134_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__or2_1
XFILLER_59_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12850_ sha256cu.m_pad_pars.block_512\[29\]\[2\] _06407_ VGND VGND VPWR VPWR _06410_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11801_ sha256cu.msg_scheduler.mreg_1\[27\] _05624_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__xnor2_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12781_ _06373_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__clkbuf_1
X_14520_ clknet_leaf_120_clk _01034_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ sha256cu.msg_scheduler.mreg_14\[25\] _05558_ VGND VGND VPWR VPWR _05559_
+ sky130_fd_sc_hd__xnor2_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _05490_ _05491_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__nand2_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ clknet_leaf_6_clk _00965_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10614_ sha256cu.msg_scheduler.mreg_10\[10\] _04574_ VGND VGND VPWR VPWR _04587_
+ sky130_fd_sc_hd__or2_1
X_14382_ clknet_leaf_108_clk _00896_ VGND VGND VPWR VPWR sha256cu.iter_processing.padding_done
+ sky130_fd_sc_hd__dfxtp_4
X_13402_ _06702_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_1
X_11594_ _03288_ _02009_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__and2_1
XFILLER_6_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13333_ _06666_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_1
X_10545_ _01566_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10476_ sha256cu.msg_scheduler.mreg_8\[15\] _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__or2_1
XFILLER_6_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13264_ _06630_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
X_12215_ _06019_ _06020_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__or2_1
X_13195_ sha256cu.m_pad_pars.block_512\[49\]\[3\] _06590_ VGND VGND VPWR VPWR _06594_
+ sky130_fd_sc_hd__and2_1
X_12146_ _05954_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__nor2_1
XFILLER_111_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12077_ _05775_ _05887_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__a21bo_1
XFILLER_38_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11028_ sha256cu.m_pad_pars.block_512\[11\]\[5\] _04790_ _04831_ sha256cu.m_pad_pars.block_512\[19\]\[5\]
+ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__a22o_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12979_ _06478_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14718_ clknet_leaf_123_clk _01232_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14649_ clknet_leaf_123_clk _01163_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_38 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _01554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _02747_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__inv_2
XANTENNA_27 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_49 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07121_ _01640_ _01594_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__nor2_1
XFILLER_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_121_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_121_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07052_ _01667_ _01614_ _01584_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07954_ sha256cu.m_out_digest.h_in\[15\] _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__xnor2_2
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07885_ _02455_ _02457_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__nor2_1
XFILLER_68_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06905_ _01596_ _01597_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__or2_2
XFILLER_95_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09624_ sha256cu.m_out_digest.g_in\[24\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[24\]
+ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__o22a_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06836_ net113 net116 net115 net118 VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__or4_1
XFILLER_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09555_ _02220_ _04023_ _04024_ _04025_ _01984_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__o311a_1
X_09486_ sha256cu.m_out_digest.h_in\[29\] sha256cu.m_out_digest.d_in\[29\] VGND VGND
+ VPWR VPWR _03959_ sky130_fd_sc_hd__or2_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08506_ _03106_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__inv_2
X_08437_ _03016_ _03018_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__nor2_1
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08368_ _02970_ _02971_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07319_ _01961_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_112_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_16
X_08299_ sha256cu.iter_processing.w\[24\] _02904_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__xor2_1
XFILLER_20_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10330_ sha256cu.msg_scheduler.mreg_6\[16\] _04415_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__or2_1
XFILLER_125_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10261_ sha256cu.msg_scheduler.mreg_5\[19\] _04374_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__or2_1
XFILLER_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12000_ _05814_ _05815_ _05442_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__o21a_1
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10192_ sha256cu.msg_scheduler.mreg_4\[21\] _04335_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__or2_1
X_13951_ clknet_leaf_54_clk _00497_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_87_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12902_ _06437_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__clkbuf_1
X_13882_ clknet_leaf_23_clk _00428_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12833_ sha256cu.m_pad_pars.block_512\[28\]\[2\] _06398_ VGND VGND VPWR VPWR _06401_
+ sky130_fd_sc_hd__and2_1
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _06364_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _05515_ _05529_ _05542_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__and3_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ clknet_leaf_13_clk _01017_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _06327_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11646_ sha256cu.msg_scheduler.mreg_14\[21\] _05476_ VGND VGND VPWR VPWR _05477_
+ sky130_fd_sc_hd__xnor2_1
X_14434_ clknet_leaf_104_clk _00948_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput25 hash[121] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput14 hash[111] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
X_14365_ clknet_leaf_77_clk _00879_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput36 hash[131] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
X_11577_ _04769_ _04808_ _05282_ sha256cu.m_pad_pars.block_512\[16\]\[7\] VGND VGND
+ VPWR VPWR _05413_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_103_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_16
Xinput47 hash[141] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xinput69 hash[161] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10528_ sha256cu.msg_scheduler.mreg_8\[5\] _04526_ _04537_ _04530_ VGND VGND VPWR
+ VPWR _00721_ sky130_fd_sc_hd__o211a_1
XFILLER_109_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput58 hash[151] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
X_14296_ clknet_leaf_20_clk _00842_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13316_ _06657_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13247_ _06621_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10459_ sha256cu.msg_scheduler.mreg_8\[8\] _04494_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__or2_1
XFILLER_124_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13178_ _06584_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__clkbuf_1
X_12129_ sha256cu.data_in_padd\[22\] _05667_ _05939_ _05445_ VGND VGND VPWR VPWR _05940_
+ sky130_fd_sc_hd__a211o_1
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07670_ sha256cu.m_out_digest.a_in\[7\] _02070_ _02114_ _02292_ VGND VGND VPWR VPWR
+ _00102_ sky130_fd_sc_hd__a22o_1
XFILLER_65_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09340_ _03816_ _03817_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__or2_1
X_09271_ _03725_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__inv_2
XFILLER_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08222_ _02784_ _02785_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__and2b_1
XFILLER_147_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08153_ _02621_ _02661_ _02762_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__or3b_1
X_08084_ _02661_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__inv_2
X_07104_ _01622_ _01687_ _01694_ _01652_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__o31ai_1
X_07035_ _01679_ _01713_ _01718_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__o21a_1
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08986_ sha256cu.m_out_digest.h_in\[12\] sha256cu.m_out_digest.d_in\[12\] VGND VGND
+ VPWR VPWR _03476_ sky130_fd_sc_hd__nor2_1
XFILLER_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07937_ _02552_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07868_ sha256cu.iter_processing.w\[12\] _02447_ _02484_ VGND VGND VPWR VPWR _02485_
+ sky130_fd_sc_hd__a21o_1
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07799_ _02417_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__inv_2
X_09607_ sha256cu.m_out_digest.g_in\[11\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[11\]
+ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__o22a_1
X_06819_ _01504_ _01506_ _01511_ _01516_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__or4_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09538_ sha256cu.m_out_digest.e_in\[30\] _02629_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__and2_1
X_09469_ _03941_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__nor2_1
XFILLER_52_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ sha256cu.m_pad_pars.block_512\[60\]\[2\] _01998_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[2\]
+ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__a22o_1
XFILLER_138_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12480_ sha256cu.m_pad_pars.block_512\[7\]\[6\] _06205_ VGND VGND VPWR VPWR _06212_
+ sky130_fd_sc_hd__and2_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11431_ sha256cu.data_in_padd\[23\] _04840_ _05274_ _04709_ VGND VGND VPWR VPWR _00886_
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14150_ clknet_leaf_34_clk _00696_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11362_ sha256cu.m_pad_pars.block_512\[41\]\[4\] _05132_ _05144_ sha256cu.m_pad_pars.block_512\[9\]\[4\]
+ _05208_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__a221o_1
XFILLER_153_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10313_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__clkbuf_2
XFILLER_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13101_ _06543_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__clkbuf_1
X_14081_ clknet_leaf_37_clk _00627_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11293_ _04769_ _05130_ _05139_ _05127_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__o211a_2
X_10244_ sha256cu.msg_scheduler.mreg_4\[11\] _04367_ _04375_ _04370_ VGND VGND VPWR
+ VPWR _00599_ sky130_fd_sc_hd__o211a_1
XFILLER_112_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13032_ _06506_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__clkbuf_1
X_10175_ sha256cu.msg_scheduler.mreg_3\[13\] _04328_ _04336_ _04331_ VGND VGND VPWR
+ VPWR _00569_ sky130_fd_sc_hd__o211a_1
XFILLER_133_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13934_ clknet_leaf_50_clk _00480_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_13865_ clknet_leaf_21_clk _00411_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12816_ sha256cu.m_pad_pars.block_512\[27\]\[2\] _06389_ VGND VGND VPWR VPWR _06392_
+ sky130_fd_sc_hd__and2_1
XFILLER_90_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13796_ clknet_leaf_85_clk _00342_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12747_ _06355_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _06318_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__clkbuf_1
X_11629_ _05444_ _05459_ _05432_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__a21o_1
X_14417_ clknet_leaf_107_clk _00931_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_512_block\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14348_ clknet_leaf_108_clk _00862_ VGND VGND VPWR VPWR sha256cu.flag_0_15 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14279_ clknet_leaf_23_clk _00825_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _03333_ _03335_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__nand2_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _02126_ _03245_ _03246_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__a21boi_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07722_ sha256cu.m_out_digest.e_in\[15\] sha256cu.m_out_digest.e_in\[2\] VGND VGND
+ VPWR VPWR _02343_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07653_ sha256cu.m_out_digest.h_in\[7\] _02275_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__xnor2_2
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07584_ _02206_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09323_ _03762_ _03769_ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__o21a_1
XFILLER_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09254_ _03732_ _03733_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__and2_1
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09185_ sha256cu.m_out_digest.e_in\[18\] _02040_ _03668_ _02068_ VGND VGND VPWR VPWR
+ _00241_ sky130_fd_sc_hd__a211o_1
X_08205_ _02777_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__inv_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08136_ sha256cu.m_out_digest.e_in\[26\] sha256cu.m_out_digest.e_in\[13\] VGND VGND
+ VPWR VPWR _02746_ sky130_fd_sc_hd__xnor2_2
XFILLER_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08067_ sha256cu.m_out_digest.h_in\[18\] _02678_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07018_ _01601_ _01588_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__nor2_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput204 hash[52] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput226 hash[72] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_2
Xinput215 hash[62] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
X_08969_ _03458_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__nand2_1
XFILLER_124_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput248 hash[92] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput237 hash[82] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_2
X_11980_ sha256cu.data_in_padd\[16\] _05433_ _05795_ _05796_ _04046_ VGND VGND VPWR
+ VPWR _05797_ sky130_fd_sc_hd__a221o_1
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10931_ _04735_ sha256cu.m_pad_pars.add_out3\[4\] VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__nor2_1
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13650_ clknet_leaf_60_clk _00196_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10862_ _01975_ _04732_ _04733_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__and3_1
XFILLER_140_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ sha256cu.msg_scheduler.mreg_11\[23\] _04685_ _04687_ _04688_ VGND VGND VPWR
+ VPWR _00835_ sky130_fd_sc_hd__o211a_1
X_13581_ clknet_leaf_74_clk _00127_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12601_ _06277_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ _06239_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12463_ sha256cu.m_pad_pars.block_512\[6\]\[6\] _06196_ VGND VGND VPWR VPWR _06203_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14202_ clknet_leaf_19_clk _00748_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11414_ _04933_ _05248_ _05257_ sha256cu.m_pad_pars.block_512\[13\]\[7\] VGND VGND
+ VPWR VPWR _05258_ sky130_fd_sc_hd__o22a_1
XFILLER_125_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12394_ _06166_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__clkbuf_1
X_14133_ clknet_leaf_34_clk _00679_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11345_ sha256cu.m_pad_pars.block_512\[25\]\[3\] _05140_ _05138_ sha256cu.m_pad_pars.block_512\[17\]\[3\]
+ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__a22o_1
XFILLER_152_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14064_ clknet_leaf_38_clk _00610_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11276_ sha256cu.m_pad_pars.add_out1\[5\] sha256cu.m_pad_pars.add_out1\[4\] VGND
+ VGND VPWR VPWR _05127_ sky130_fd_sc_hd__nor2_2
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10227_ sha256cu.msg_scheduler.mreg_4\[4\] _04354_ _04365_ _04357_ VGND VGND VPWR
+ VPWR _00592_ sky130_fd_sc_hd__o211a_1
X_13015_ _06497_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__clkbuf_1
X_10158_ sha256cu.msg_scheduler.mreg_3\[6\] _04315_ _04326_ _04318_ VGND VGND VPWR
+ VPWR _00562_ sky130_fd_sc_hd__o211a_1
XFILLER_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10089_ sha256cu.msg_scheduler.mreg_3\[9\] _04282_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__or2_1
XFILLER_94_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13917_ clknet_leaf_45_clk _00463_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14897_ clknet_leaf_0_clk _01411_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13848_ clknet_leaf_21_clk _00394_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13779_ clknet_leaf_60_clk _00325_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09941_ sha256cu.msg_scheduler.mreg_1\[9\] _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__or2_1
XFILLER_89_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09872_ sha256cu.msg_scheduler.mreg_13\[21\] _04160_ VGND VGND VPWR VPWR _04161_
+ sky130_fd_sc_hd__or2_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08823_ sha256cu.iter_processing.w\[6\] _02224_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__and2_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _03225_ _03231_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__o21a_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _02260_ _02289_ _02249_ _02251_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__a211o_1
XFILLER_66_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_309 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08685_ sha256cu.m_out_digest.d_in\[27\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[27\]
+ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__a22o_1
XFILLER_54_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_26_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07636_ _02245_ _02247_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__nor2_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07567_ _02188_ _02189_ _02190_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__a21o_1
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09306_ _03774_ _03775_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__nand2_1
XFILLER_22_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07498_ sha256cu.m_out_digest.e_in\[14\] sha256cu.m_out_digest.e_in\[9\] VGND VGND
+ VPWR VPWR _02125_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09237_ _03717_ _03718_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__and2_1
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09168_ _03650_ _03651_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__nor2_1
X_09099_ sha256cu.m_out_digest.h_in\[16\] sha256cu.m_out_digest.d_in\[16\] VGND VGND
+ VPWR VPWR _03585_ sky130_fd_sc_hd__or2_1
X_08119_ _02695_ _02698_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__o21ba_1
XFILLER_150_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11130_ _04987_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__nor2_4
XFILLER_1_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11061_ _04764_ _04798_ _04920_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__and3_1
X_10012_ sha256cu.msg_scheduler.mreg_2\[8\] _04241_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__or2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14820_ clknet_leaf_101_clk _01334_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11963_ sha256cu.msg_scheduler.mreg_1\[23\] _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14751_ clknet_leaf_106_clk _01265_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[41\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11894_ sha256cu.msg_scheduler.mreg_1\[20\] sha256cu.msg_scheduler.mreg_1\[16\] VGND
+ VGND VPWR VPWR _05714_ sky130_fd_sc_hd__xnor2_1
X_13702_ clknet_leaf_83_clk _00248_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[25\]
+ sky130_fd_sc_hd__dfxtp_4
X_10914_ _04730_ _04766_ _04778_ _04780_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__and4b_2
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14682_ clknet_leaf_120_clk _01196_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13633_ clknet_leaf_85_clk _00179_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10845_ sha256cu.m_pad_pars.add_out2\[4\] VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__clkbuf_2
XFILLER_60_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13564_ clknet_leaf_64_clk _00110_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10776_ sha256cu.msg_scheduler.mreg_11\[16\] _04672_ _04678_ _04675_ VGND VGND VPWR
+ VPWR _00828_ sky130_fd_sc_hd__o211a_1
XFILLER_9_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12515_ _06230_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13495_ sha256cu.K\[24\] _06713_ _06718_ _00052_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__a22o_1
XFILLER_126_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12446_ sha256cu.m_pad_pars.block_512\[5\]\[6\] _06187_ VGND VGND VPWR VPWR _06194_
+ sky130_fd_sc_hd__and2_1
X_12377_ sha256cu.m_pad_pars.block_512\[1\]\[5\] _06152_ VGND VGND VPWR VPWR _06158_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14116_ clknet_leaf_37_clk _00662_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11328_ sha256cu.m_pad_pars.block_512\[25\]\[1\] _05140_ _05158_ sha256cu.m_pad_pars.block_512\[21\]\[1\]
+ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__a221o_1
XFILLER_125_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14047_ clknet_leaf_39_clk _00593_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11259_ sha256cu.m_pad_pars.block_512\[22\]\[7\] _05011_ _05012_ VGND VGND VPWR VPWR
+ _05111_ sky130_fd_sc_hd__o21ba_1
XFILLER_67_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_75_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14949_ clknet_leaf_91_clk _01463_ VGND VGND VPWR VPWR sha256cu.K\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08470_ _03070_ _03033_ _03034_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__and3_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07421_ sha256cu.m_out_digest.e_in\[12\] sha256cu.m_out_digest.e_in\[7\] VGND VGND
+ VPWR VPWR _02050_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07352_ sha256cu.m_pad_pars.add_out0\[3\] sha256cu.m_pad_pars.add_out0\[2\] VGND
+ VGND VPWR VPWR _01991_ sky130_fd_sc_hd__nand2_1
XFILLER_148_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07283_ sha256cu.m_pad_pars.m_size\[5\] sha256cu.m_pad_pars.block_512\[63\]\[5\]
+ _01928_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__mux2_1
X_09022_ _02450_ _03478_ _03477_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__a21oi_1
X_09924_ sha256cu.msg_scheduler.mreg_1\[2\] _04174_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__or2_1
XFILLER_98_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09855_ sha256cu.msg_scheduler.mreg_13\[14\] _04147_ VGND VGND VPWR VPWR _04151_
+ sky130_fd_sc_hd__or2_1
XFILLER_58_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _03270_ _03275_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__o21a_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09786_ sha256cu.msg_scheduler.mreg_14\[17\] _04106_ VGND VGND VPWR VPWR _04111_
+ sky130_fd_sc_hd__or2_1
XFILLER_58_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06998_ _00452_ _01658_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__nand2_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
X_08737_ _03220_ _03218_ _03236_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__a21oi_2
XANTENNA_106 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08668_ sha256cu.m_out_digest.d_in\[12\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[12\]
+ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__o22a_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07619_ _02194_ _02205_ _02242_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__o21ba_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08599_ _02113_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__buf_6
X_10630_ sha256cu.msg_scheduler.mreg_10\[17\] _04588_ VGND VGND VPWR VPWR _04596_
+ sky130_fd_sc_hd__or2_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10561_ _04529_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__buf_2
X_10492_ sha256cu.msg_scheduler.mreg_8\[22\] _04507_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__or2_1
XFILLER_127_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12300_ _06101_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__xor2_1
X_13280_ sha256cu.m_pad_pars.block_512\[54\]\[3\] _06635_ VGND VGND VPWR VPWR _06639_
+ sky130_fd_sc_hd__and2_1
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12231_ sha256cu.msg_scheduler.mreg_1\[30\] _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xpassword_cracker_271 VGND VGND VPWR VPWR password_cracker_271/HI password_count[11]
+ sky130_fd_sc_hd__conb_1
Xpassword_cracker_260 VGND VGND VPWR VPWR password_cracker_260/HI password_count[0]
+ sky130_fd_sc_hd__conb_1
Xpassword_cracker_282 VGND VGND VPWR VPWR password_cracker_282/HI password_count[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12162_ sha256cu.msg_scheduler.mreg_1\[27\] sha256cu.msg_scheduler.mreg_1\[10\] VGND
+ VGND VPWR VPWR _05971_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12093_ sha256cu.msg_scheduler.mreg_14\[8\] sha256cu.msg_scheduler.mreg_14\[6\] VGND
+ VGND VPWR VPWR _05905_ sky130_fd_sc_hd__xnor2_1
X_11113_ _04968_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__nor2_4
XFILLER_104_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11044_ _01971_ _04903_ _04904_ _04709_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__o211a_1
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_56_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_64_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12995_ sha256cu.m_pad_pars.block_512\[37\]\[6\] _06480_ VGND VGND VPWR VPWR _06487_
+ sky130_fd_sc_hd__and2_1
X_14803_ clknet_leaf_1_clk _01317_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11946_ _05762_ _05763_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nor2_1
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14734_ clknet_leaf_11_clk _01248_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11877_ sha256cu.msg_scheduler.mreg_14\[29\] sha256cu.msg_scheduler.mreg_14\[22\]
+ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__xnor2_1
X_14665_ clknet_leaf_13_clk _01179_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13616_ clknet_leaf_51_clk _00162_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14596_ clknet_leaf_101_clk _01110_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10828_ sha256cu.m_pad_pars.add_512_block\[3\] _04700_ _04711_ _04709_ VGND VGND
+ VPWR VPWR _00847_ sky130_fd_sc_hd__o211a_1
X_10759_ sha256cu.msg_scheduler.mreg_12\[9\] _04666_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__or2_1
X_13547_ clknet_leaf_79_clk _00093_ VGND VGND VPWR VPWR sha256cu.m_out_digest.H7\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13478_ sha256cu.K\[17\] _06726_ _06727_ _06750_ _06737_ VGND VGND VPWR VPWR _01458_
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12429_ sha256cu.m_pad_pars.block_512\[4\]\[6\] _06178_ VGND VGND VPWR VPWR _06185_
+ sky130_fd_sc_hd__and2_1
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07970_ _02555_ _02556_ _02582_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__a21oi_2
X_06921_ _01592_ _01580_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__nand2_4
X_09640_ sha256cu.m_out_digest.h_in\[6\] _04037_ _04036_ sha256cu.m_out_digest.g_in\[6\]
+ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__a22o_1
X_06852_ net24 net27 net26 net29 VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__or4_4
X_09571_ sha256cu.m_out_digest.f_in\[12\] _03559_ _04028_ sha256cu.m_out_digest.e_in\[12\]
+ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__a22o_1
X_06783_ _01477_ _01478_ _01479_ _01480_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__or4_1
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_47_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
X_08522_ sha256cu.m_out_digest.h_in\[29\] _03079_ _03121_ VGND VGND VPWR VPWR _03122_
+ sky130_fd_sc_hd__a21bo_1
X_08453_ _03049_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__nand2_1
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07404_ _02032_ _02033_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__nor2_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08384_ _02986_ _02987_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__xnor2_2
X_07335_ sha256cu.m_pad_pars.add_out1\[3\] sha256cu.m_pad_pars.add_out1\[2\] VGND
+ VGND VPWR VPWR _01977_ sky130_fd_sc_hd__and2_2
X_07266_ _01918_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__clkbuf_4
X_09005_ _03466_ _03467_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a21bo_1
X_07197_ _01623_ _01723_ _01611_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09907_ _04181_ _02007_ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__and3b_1
X_09838_ sha256cu.msg_scheduler.mreg_12\[6\] _04140_ _04141_ _04130_ VGND VGND VPWR
+ VPWR _00421_ sky130_fd_sc_hd__o211a_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09769_ sha256cu.msg_scheduler.mreg_13\[9\] _04099_ _04101_ _04090_ VGND VGND VPWR
+ VPWR _00392_ sky130_fd_sc_hd__o211a_1
XFILLER_74_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_38_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_132_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11800_ sha256cu.msg_scheduler.mreg_1\[16\] sha256cu.msg_scheduler.mreg_1\[12\] VGND
+ VGND VPWR VPWR _05624_ sky130_fd_sc_hd__xnor2_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ sha256cu.m_pad_pars.block_512\[25\]\[1\] _06371_ VGND VGND VPWR VPWR _06373_
+ sky130_fd_sc_hd__and2_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ sha256cu.msg_scheduler.mreg_14\[23\] sha256cu.msg_scheduler.mreg_14\[16\]
+ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__xnor2_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11662_ _05490_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__or2_1
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ clknet_leaf_6_clk _00964_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10613_ sha256cu.msg_scheduler.mreg_9\[9\] _04581_ _04586_ _04584_ VGND VGND VPWR
+ VPWR _00757_ sky130_fd_sc_hd__o211a_1
X_11593_ sha256cu.data_in_padd\[31\] _01980_ _01987_ _05428_ VGND VGND VPWR VPWR _00894_
+ sky130_fd_sc_hd__a22o_1
X_14381_ clknet_leaf_79_clk _00895_ VGND VGND VPWR VPWR sha256cu.hashing_done sky130_fd_sc_hd__dfxtp_1
X_13401_ sha256cu.m_pad_pars.block_512\[61\]\[5\] _06693_ VGND VGND VPWR VPWR _06702_
+ sky130_fd_sc_hd__and2_1
XFILLER_128_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10544_ sha256cu.msg_scheduler.mreg_8\[12\] _04540_ _04546_ _04543_ VGND VGND VPWR
+ VPWR _00728_ sky130_fd_sc_hd__o211a_1
X_13332_ sha256cu.m_pad_pars.block_512\[57\]\[4\] _06660_ VGND VGND VPWR VPWR _06666_
+ sky130_fd_sc_hd__and2_1
XFILLER_10_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10475_ _04414_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__clkbuf_2
XFILLER_124_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13263_ sha256cu.m_pad_pars.block_512\[53\]\[3\] _06626_ VGND VGND VPWR VPWR _06630_
+ sky130_fd_sc_hd__and2_1
XFILLER_136_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12214_ _06019_ _06020_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__nand2_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13194_ _06593_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12145_ _05923_ _05927_ _05952_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__a21oi_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12076_ _05859_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__and2_1
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11027_ sha256cu.m_pad_pars.block_512\[23\]\[5\] _04828_ _04818_ sha256cu.m_pad_pars.block_512\[35\]\[5\]
+ _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__a221o_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_64_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12978_ sha256cu.m_pad_pars.block_512\[36\]\[6\] _06471_ VGND VGND VPWR VPWR _06478_
+ sky130_fd_sc_hd__and2_1
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ _05745_ _05746_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__nand2_1
X_14717_ clknet_leaf_121_clk _01231_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14648_ clknet_leaf_122_clk _01162_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_39 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _01554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14579_ clknet_leaf_5_clk _01093_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07120_ _01617_ _01727_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__nand2_1
XFILLER_146_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07051_ _01607_ _01606_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__or2_1
XFILLER_126_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07953_ _02232_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__xnor2_2
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07884_ _02490_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__xor2_1
XFILLER_95_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06904_ _01593_ _01589_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__nor2_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09623_ sha256cu.m_out_digest.g_in\[23\] _04035_ _04034_ sha256cu.m_out_digest.f_in\[23\]
+ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__o22a_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06835_ net117 net120 net119 net122 VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__or4_1
XFILLER_28_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09554_ sha256cu.m_out_digest.e_in\[31\] _02439_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__or2_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09485_ sha256cu.m_out_digest.h_in\[29\] sha256cu.m_out_digest.d_in\[29\] VGND VGND
+ VPWR VPWR _03958_ sky130_fd_sc_hd__nand2_1
XFILLER_64_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08505_ _03064_ _03074_ _03104_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__and3_1
X_08436_ _03011_ _03012_ _03015_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__and3_1
X_08367_ sha256cu.m_out_digest.g_in\[26\] sha256cu.m_out_digest.f_in\[26\] sha256cu.m_out_digest.e_in\[26\]
+ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__mux2_2
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07318_ sha256cu.m_pad_pars.add_out1\[2\] _01961_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__and2_1
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08298_ _02902_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07249_ state\[2\] _00032_ _01563_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__or3_1
X_10260_ sha256cu.msg_scheduler.mreg_4\[18\] _04380_ _04384_ _04383_ VGND VGND VPWR
+ VPWR _00606_ sky130_fd_sc_hd__o211a_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10191_ sha256cu.msg_scheduler.mreg_3\[20\] _04341_ _04345_ _04344_ VGND VGND VPWR
+ VPWR _00576_ sky130_fd_sc_hd__o211a_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13950_ clknet_leaf_54_clk _00496_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12901_ sha256cu.m_pad_pars.block_512\[32\]\[2\] _06434_ VGND VGND VPWR VPWR _06437_
+ sky130_fd_sc_hd__and2_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13881_ clknet_leaf_23_clk _00427_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _06400_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__clkbuf_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ sha256cu.m_pad_pars.block_512\[24\]\[1\] _06362_ VGND VGND VPWR VPWR _06364_
+ sky130_fd_sc_hd__and2_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _05539_ _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__xnor2_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ clknet_leaf_107_clk _01016_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ sha256cu.m_pad_pars.block_512\[20\]\[1\] _06325_ VGND VGND VPWR VPWR _06327_
+ sky130_fd_sc_hd__and2_1
X_14433_ clknet_leaf_103_clk _00947_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11645_ sha256cu.msg_scheduler.mreg_14\[19\] sha256cu.msg_scheduler.mreg_14\[12\]
+ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__xnor2_1
Xinput15 hash[112] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 hash[122] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput37 hash[132] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14364_ clknet_leaf_109_clk _00878_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11576_ _01936_ _05293_ _05411_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__and3_1
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10527_ sha256cu.msg_scheduler.mreg_9\[5\] _04534_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__or2_1
X_14295_ clknet_leaf_20_clk _00841_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput48 hash[142] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13315_ sha256cu.m_pad_pars.block_512\[56\]\[4\] _01924_ VGND VGND VPWR VPWR _06657_
+ sky130_fd_sc_hd__and2_1
Xinput59 hash[152] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
XFILLER_143_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10458_ sha256cu.msg_scheduler.mreg_7\[7\] _04487_ _04497_ _04490_ VGND VGND VPWR
+ VPWR _00691_ sky130_fd_sc_hd__o211a_1
XFILLER_115_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13246_ sha256cu.m_pad_pars.block_512\[52\]\[3\] _06617_ VGND VGND VPWR VPWR _06621_
+ sky130_fd_sc_hd__and2_1
XFILLER_108_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10389_ sha256cu.msg_scheduler.mreg_6\[9\] _04448_ _04458_ _04451_ VGND VGND VPWR
+ VPWR _00661_ sky130_fd_sc_hd__o211a_1
X_13177_ sha256cu.m_pad_pars.block_512\[48\]\[3\] _06580_ VGND VGND VPWR VPWR _06584_
+ sky130_fd_sc_hd__and2_1
XFILLER_111_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12128_ _05465_ _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__nor2_1
X_12059_ _05869_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__xor2_1
XFILLER_111_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09270_ _03749_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__and2b_1
XFILLER_21_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08221_ _02827_ _02828_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__or2_1
XFILLER_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08152_ _02695_ _02728_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__and2b_1
XFILLER_147_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08083_ _02692_ _02694_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_9_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
X_07103_ _01648_ _01639_ _01634_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__and3_1
X_07034_ _00456_ _01716_ _01717_ _01661_ _01571_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__a221o_1
XFILLER_127_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08985_ _03455_ _03456_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07936_ _02002_ _02551_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__or2_1
XFILLER_69_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07867_ _02445_ _02446_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__and2b_1
XFILLER_84_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09606_ sha256cu.m_out_digest.g_in\[10\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[10\]
+ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__a22o_1
X_07798_ sha256cu.m_out_digest.e_in\[22\] _02416_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__xnor2_2
X_06818_ _01512_ _01513_ _01514_ _01515_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__or4_1
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09537_ _04006_ _04008_ _02069_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09468_ _03936_ _03940_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__and2_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09399_ _03873_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__or2_1
X_08419_ _03019_ _03021_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11430_ _05254_ _05263_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__or3_1
XFILLER_125_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11361_ sha256cu.m_pad_pars.block_512\[25\]\[4\] _05140_ _05141_ sha256cu.m_pad_pars.block_512\[29\]\[4\]
+ _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a221o_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10312_ _01566_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__clkbuf_4
X_13100_ sha256cu.m_pad_pars.block_512\[43\]\[7\] _04914_ _06542_ VGND VGND VPWR VPWR
+ _06543_ sky130_fd_sc_hd__mux2_1
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14080_ clknet_leaf_36_clk _00626_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11292_ sha256cu.m_pad_pars.block_512\[1\]\[0\] _05135_ _05138_ sha256cu.m_pad_pars.block_512\[17\]\[0\]
+ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__a221o_1
X_10243_ sha256cu.msg_scheduler.mreg_5\[11\] _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__or2_1
XFILLER_105_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13031_ sha256cu.m_pad_pars.block_512\[39\]\[7\] _04936_ _06442_ VGND VGND VPWR VPWR
+ _06506_ sky130_fd_sc_hd__mux2_1
X_10174_ sha256cu.msg_scheduler.mreg_4\[13\] _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__or2_1
XFILLER_105_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13933_ clknet_leaf_50_clk _00479_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13864_ clknet_leaf_22_clk _00410_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12815_ _06391_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_1
X_13795_ clknet_leaf_85_clk _00341_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ sha256cu.m_pad_pars.block_512\[23\]\[1\] _06353_ VGND VGND VPWR VPWR _06355_
+ sky130_fd_sc_hd__and2_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ sha256cu.m_pad_pars.block_512\[19\]\[1\] _06316_ VGND VGND VPWR VPWR _06318_
+ sky130_fd_sc_hd__and2_1
X_11628_ _05444_ _05459_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__nor2_1
X_14416_ clknet_leaf_107_clk _00930_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_512_block\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14347_ clknet_leaf_108_clk _00861_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11559_ _04807_ _05233_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__nor2_1
XFILLER_144_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14278_ clknet_leaf_23_clk _00824_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13229_ sha256cu.m_pad_pars.block_512\[51\]\[3\] _06608_ VGND VGND VPWR VPWR _06612_
+ sky130_fd_sc_hd__and2_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _02159_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__xor2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07721_ sha256cu.iter_processing.w\[9\] _02341_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07652_ _02272_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__xnor2_4
XFILLER_65_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07583_ _02157_ _02169_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__o21ba_1
X_09322_ _03799_ _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__nor2_1
XFILLER_139_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09253_ _03732_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__nor2_1
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09184_ _02069_ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__nor2_1
X_08204_ _02809_ _02811_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08135_ sha256cu.m_out_digest.h_in\[20\] _02744_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__xnor2_2
XFILLER_147_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08066_ sha256cu.m_out_digest.a_in\[31\] _02677_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__xnor2_2
X_07017_ _01626_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__inv_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput227 hash[73] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_4
Xinput216 hash[63] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput205 hash[53] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
X_08968_ sha256cu.iter_processing.w\[11\] _02413_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__nand2_1
XFILLER_102_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput249 hash[93] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
Xinput238 hash[83] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
X_08899_ sha256cu.m_out_digest.e_in\[8\] _02440_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__or2_1
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07919_ _02497_ _02499_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__nor2_1
XFILLER_57_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10930_ _04796_ _04791_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__or2_1
XFILLER_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12600_ sha256cu.m_pad_pars.block_512\[14\]\[5\] _06271_ VGND VGND VPWR VPWR _06277_
+ sky130_fd_sc_hd__and2_1
X_10861_ sha256cu.m_pad_pars.add_out3\[4\] _04731_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__nand2_1
XFILLER_32_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13580_ clknet_leaf_78_clk _00126_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[31\]
+ sky130_fd_sc_hd__dfxtp_4
X_10792_ _01994_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__clkbuf_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ sha256cu.m_pad_pars.block_512\[10\]\[6\] _06232_ VGND VGND VPWR VPWR _06239_
+ sky130_fd_sc_hd__and2_1
XFILLER_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12462_ _06202_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__clkbuf_1
X_14201_ clknet_leaf_28_clk _00747_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11413_ _04702_ _05096_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__nor2_1
XFILLER_8_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12393_ sha256cu.m_pad_pars.block_512\[2\]\[5\] _06160_ VGND VGND VPWR VPWR _06166_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14132_ clknet_leaf_34_clk _00678_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11344_ sha256cu.m_pad_pars.block_512\[33\]\[3\] _05147_ _05191_ VGND VGND VPWR VPWR
+ _05192_ sky130_fd_sc_hd__a21o_1
XFILLER_153_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14063_ clknet_leaf_39_clk _00609_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11275_ _04913_ _05124_ _05125_ _01977_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__o211a_2
XFILLER_152_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10226_ sha256cu.msg_scheduler.mreg_5\[4\] _04361_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__or2_1
X_13014_ sha256cu.m_pad_pars.block_512\[38\]\[7\] _05085_ _06442_ VGND VGND VPWR VPWR
+ _06497_ sky130_fd_sc_hd__mux2_1
XFILLER_95_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10157_ sha256cu.msg_scheduler.mreg_4\[6\] _04322_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__or2_1
XFILLER_121_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10088_ sha256cu.msg_scheduler.mreg_2\[8\] _04274_ _04286_ _04277_ VGND VGND VPWR
+ VPWR _00532_ sky130_fd_sc_hd__o211a_1
XFILLER_82_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13916_ clknet_leaf_45_clk _00462_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14896_ clknet_leaf_0_clk _01410_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13847_ clknet_leaf_21_clk _00393_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13778_ clknet_leaf_60_clk _00324_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12729_ _06345_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09940_ _04133_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__buf_2
XFILLER_116_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09871_ _04133_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__clkbuf_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ sha256cu.iter_processing.w\[6\] _02224_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__nor2_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _03229_ _03230_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__or2_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07704_ _02254_ _02252_ _02253_ _02290_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__nor4_2
XFILLER_72_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08684_ sha256cu.m_out_digest.d_in\[26\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[26\]
+ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__o22a_1
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07635_ sha256cu.m_out_digest.a_in\[6\] _02220_ _02256_ _02257_ _02258_ VGND VGND
+ VPWR VPWR _00101_ sky130_fd_sc_hd__a221o_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07566_ _02188_ _02189_ _02190_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__and3_1
XFILLER_139_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09305_ _02113_ _03783_ _03784_ _02332_ sha256cu.m_out_digest.e_in\[22\] VGND VGND
+ VPWR VPWR _00245_ sky130_fd_sc_hd__a32o_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07497_ sha256cu.iter_processing.w\[3\] _02123_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__xnor2_1
X_09236_ _03715_ _03716_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__or2_1
XFILLER_22_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09167_ sha256cu.iter_processing.w\[18\] _02671_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__and2_1
XFILLER_135_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09098_ sha256cu.m_out_digest.e_in\[15\] _03559_ _03192_ _03584_ VGND VGND VPWR VPWR
+ _00238_ sky130_fd_sc_hd__a22o_1
X_08118_ _02692_ _02694_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__and2b_1
XFILLER_123_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08049_ _02619_ _02630_ _02661_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__o21ai_1
XFILLER_150_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11060_ _04758_ _04913_ _04816_ sha256cu.m_pad_pars.block_512\[35\]\[7\] VGND VGND
+ VPWR VPWR _04920_ sky130_fd_sc_hd__o22a_1
XFILLER_1_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10011_ sha256cu.msg_scheduler.mreg_1\[7\] _04234_ _04242_ _04237_ VGND VGND VPWR
+ VPWR _00499_ sky130_fd_sc_hd__o211a_1
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14750_ clknet_leaf_123_clk _01264_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11962_ sha256cu.msg_scheduler.mreg_1\[19\] sha256cu.msg_scheduler.mreg_1\[2\] VGND
+ VGND VPWR VPWR _05779_ sky130_fd_sc_hd__xnor2_1
X_13701_ clknet_leaf_83_clk _00247_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[24\]
+ sky130_fd_sc_hd__dfxtp_4
X_11893_ _05711_ _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__nand2_1
X_10913_ _04768_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__or2_1
X_14681_ clknet_leaf_121_clk _01195_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13632_ clknet_leaf_84_clk _00178_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10844_ sha256cu.m_pad_pars.add_out2\[3\] _04718_ _04720_ _01971_ _01974_ VGND VGND
+ VPWR VPWR _00854_ sky130_fd_sc_hd__o221a_1
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13563_ clknet_leaf_65_clk _00109_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[14\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_13_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10775_ sha256cu.msg_scheduler.mreg_12\[16\] _04666_ VGND VGND VPWR VPWR _04678_
+ sky130_fd_sc_hd__or2_1
X_12514_ sha256cu.m_pad_pars.block_512\[9\]\[6\] _06223_ VGND VGND VPWR VPWR _06230_
+ sky130_fd_sc_hd__and2_1
XFILLER_9_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13494_ sha256cu.K\[23\] _06716_ _06717_ _06760_ _06737_ VGND VGND VPWR VPWR _01464_
+ sky130_fd_sc_hd__o221a_1
X_12445_ _06193_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__clkbuf_1
X_12376_ _06157_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ clknet_leaf_37_clk _00661_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11327_ sha256cu.m_pad_pars.block_512\[5\]\[1\] _05160_ _05165_ sha256cu.m_pad_pars.block_512\[37\]\[1\]
+ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__a221o_1
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14046_ clknet_leaf_39_clk _00592_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11258_ _04725_ _04721_ _04990_ _05109_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__and4_1
X_10209_ sha256cu.msg_scheduler.mreg_3\[28\] _04354_ _04355_ _04344_ VGND VGND VPWR
+ VPWR _00584_ sky130_fd_sc_hd__o211a_1
XFILLER_122_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11189_ sha256cu.m_pad_pars.block_512\[26\]\[3\] _04964_ _05014_ sha256cu.m_pad_pars.block_512\[18\]\[3\]
+ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__a22o_1
XFILLER_67_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14948_ clknet_leaf_91_clk _01462_ VGND VGND VPWR VPWR sha256cu.K\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14879_ clknet_leaf_100_clk _01393_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[57\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07420_ sha256cu.iter_processing.w\[1\] _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07351_ _01989_ _01990_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__nor2_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07282_ _01930_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09021_ _02492_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09923_ sha256cu.msg_scheduler.mreg_0\[1\] _04167_ _04192_ _04171_ VGND VGND VPWR
+ VPWR _00461_ sky130_fd_sc_hd__o211a_1
X_09854_ sha256cu.msg_scheduler.mreg_12\[13\] _04140_ _04150_ _04144_ VGND VGND VPWR
+ VPWR _00428_ sky130_fd_sc_hd__o211a_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _03268_ _03269_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__or2_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ sha256cu.msg_scheduler.mreg_13\[16\] _04099_ _04110_ _04103_ VGND VGND VPWR
+ VPWR _00399_ sky130_fd_sc_hd__o211a_1
X_06997_ _00455_ _01681_ _01682_ _00452_ _01621_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__a221o_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _03221_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_107 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ sha256cu.m_out_digest.d_in\[11\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[11\]
+ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__a22o_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07618_ _02202_ _02204_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__nor2_1
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08598_ sha256cu.m_out_digest.b_in\[18\] _03177_ _03176_ _02198_ VGND VGND VPWR VPWR
+ _00145_ sky130_fd_sc_hd__o22a_1
X_07549_ _02138_ _02136_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__and2b_1
XFILLER_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10560_ sha256cu.msg_scheduler.mreg_9\[19\] _04548_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__or2_1
XFILLER_10_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10491_ sha256cu.msg_scheduler.mreg_7\[21\] _04513_ _04515_ _04516_ VGND VGND VPWR
+ VPWR _00705_ sky130_fd_sc_hd__o211a_1
X_09219_ _03699_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nor2_1
XFILLER_135_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12230_ sha256cu.msg_scheduler.mreg_1\[13\] sha256cu.msg_scheduler.mreg_1\[2\] VGND
+ VGND VPWR VPWR _06036_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpassword_cracker_261 VGND VGND VPWR VPWR password_cracker_261/HI password_count[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_146_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12161_ _05968_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__nand2_1
Xpassword_cracker_272 VGND VGND VPWR VPWR password_cracker_272/HI password_count[12]
+ sky130_fd_sc_hd__conb_1
Xpassword_cracker_283 VGND VGND VPWR VPWR password_cracker_283/HI password_count[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_146_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12092_ _05902_ _05903_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__nor2_1
X_11112_ _04791_ _04969_ _04970_ _04698_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_150_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11043_ sha256cu.data_in_padd\[6\] _01961_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__or2_1
XFILLER_1_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_14802_ clknet_leaf_2_clk _01316_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12994_ _06486_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__clkbuf_1
X_11945_ _05760_ _05761_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__and2_1
X_14733_ clknet_leaf_7_clk _01247_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14664_ clknet_leaf_13_clk _01178_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13615_ clknet_leaf_73_clk _00161_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11876_ _05695_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__and2_1
XFILLER_41_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14595_ clknet_leaf_104_clk _01109_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10827_ sha256cu.m_pad_pars.m_size\[6\] _04706_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__or2_1
X_10758_ sha256cu.msg_scheduler.mreg_11\[8\] _04659_ _04668_ _04662_ VGND VGND VPWR
+ VPWR _00820_ sky130_fd_sc_hd__o211a_1
X_13546_ clknet_leaf_105_clk _00092_ VGND VGND VPWR VPWR sha256cu.m_out_digest.temp_delay
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13477_ _04188_ _00044_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__and2b_1
X_10689_ sha256cu.msg_scheduler.mreg_10\[10\] _04620_ _04629_ _04623_ VGND VGND VPWR
+ VPWR _00790_ sky130_fd_sc_hd__o211a_1
X_12428_ _06184_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12359_ sha256cu.m_pad_pars.block_512\[0\]\[4\] _06144_ VGND VGND VPWR VPWR _06149_
+ sky130_fd_sc_hd__and2_1
XFILLER_4_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14029_ clknet_leaf_56_clk _00575_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06920_ _00454_ _01600_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__nor2_2
XFILLER_68_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06851_ net28 net31 net30 net33 VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__or4_2
XFILLER_28_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06782_ net123 net156 net145 net174 VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__or4_2
X_09570_ _02112_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__clkbuf_4
XFILLER_95_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08521_ _03080_ _03082_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__or2b_1
XFILLER_24_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08452_ sha256cu.iter_processing.w\[28\] _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__xor2_1
XFILLER_23_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07403_ _02022_ _02031_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__and2_1
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08383_ _02948_ _02949_ _02952_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__o21ba_1
X_07334_ _01564_ _01969_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__nand2_4
XFILLER_32_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07265_ _01916_ _01917_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__or2_1
X_09004_ _03462_ _03463_ _03465_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__or3_1
X_07196_ _01665_ _01647_ _01733_ _01598_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__a31o_1
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09906_ sha256cu.msg_scheduler.counter_iteration\[2\] _04178_ sha256cu.msg_scheduler.counter_iteration\[3\]
+ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__a21o_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09837_ sha256cu.msg_scheduler.mreg_13\[6\] _04134_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__or2_1
XFILLER_86_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ sha256cu.msg_scheduler.mreg_14\[9\] _04093_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__or2_1
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ sha256cu.m_out_digest.e_in\[1\] _02220_ _03218_ _03219_ _02258_ VGND VGND
+ VPWR VPWR _00224_ sky130_fd_sc_hd__a221o_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _05555_ _05556_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__xor2_1
XFILLER_92_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09699_ sha256cu.iter_processing.w\[11\] _04054_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__or2_1
XFILLER_82_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _05469_ _05472_ _05468_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__a21boi_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10612_ sha256cu.msg_scheduler.mreg_10\[9\] _04574_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__or2_1
X_14380_ clknet_leaf_110_clk _00894_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_13400_ _06701_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__clkbuf_1
X_11592_ sha256cu.m_pad_pars.block_512\[0\]\[7\] _05386_ _05392_ _05427_ VGND VGND
+ VPWR VPWR _05428_ sky130_fd_sc_hd__o22a_1
X_10543_ sha256cu.msg_scheduler.mreg_9\[12\] _04534_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__or2_1
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13331_ _06665_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10474_ sha256cu.msg_scheduler.mreg_7\[14\] _04500_ _04506_ _04503_ VGND VGND VPWR
+ VPWR _00698_ sky130_fd_sc_hd__o211a_1
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13262_ _06629_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12213_ sha256cu.msg_scheduler.mreg_14\[13\] sha256cu.msg_scheduler.mreg_14\[11\]
+ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__xor2_1
X_13193_ sha256cu.m_pad_pars.block_512\[49\]\[2\] _06590_ VGND VGND VPWR VPWR _06593_
+ sky130_fd_sc_hd__and2_1
XFILLER_151_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12144_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__inv_2
XFILLER_151_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12075_ _05840_ _05818_ _05861_ _05858_ _05838_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__o32a_1
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11026_ sha256cu.m_pad_pars.block_512\[3\]\[5\] _04765_ _04774_ sha256cu.m_pad_pars.block_512\[7\]\[5\]
+ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__a22o_1
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12977_ _06477_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ _05745_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__or2_2
X_14716_ clknet_leaf_122_clk _01230_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11859_ _05649_ _05654_ _05680_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__and3_1
X_14647_ clknet_leaf_123_clk _01161_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[28\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_29 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14578_ clknet_leaf_4_clk _01092_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_18 _01975_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13529_ clknet_leaf_123_clk _00079_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_07050_ _01732_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07952_ _02162_ sha256cu.m_out_digest.a_in\[5\] VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07883_ _02497_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06903_ _01583_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__inv_2
X_06834_ _01528_ _01529_ _01530_ _01531_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__or4_1
X_09622_ sha256cu.m_out_digest.g_in\[22\] _04037_ _04036_ sha256cu.m_out_digest.f_in\[22\]
+ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__a22o_1
X_09553_ _04004_ _04007_ _04022_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08504_ _03064_ _03074_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__a21o_1
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ _03946_ _03947_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__nand2_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08435_ sha256cu.K\[28\] VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__inv_2
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08366_ sha256cu.m_out_digest.b_in\[26\] _02161_ _02969_ VGND VGND VPWR VPWR _02970_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07317_ _01938_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__nor2_4
XFILLER_137_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08297_ sha256cu.m_out_digest.g_in\[24\] sha256cu.m_out_digest.f_in\[24\] sha256cu.m_out_digest.e_in\[24\]
+ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__mux2_2
XFILLER_11_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07248_ _01679_ _01902_ _01903_ _01905_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__a31o_1
XFILLER_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07179_ _01650_ _01714_ _01820_ _01846_ _01663_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__o311a_1
X_10190_ sha256cu.msg_scheduler.mreg_4\[20\] _04335_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__or2_1
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13880_ clknet_leaf_22_clk _00426_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12900_ _06436_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__clkbuf_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ sha256cu.m_pad_pars.block_512\[28\]\[1\] _06398_ VGND VGND VPWR VPWR _06400_
+ sky130_fd_sc_hd__and2_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12762_ _06363_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ sha256cu.msg_scheduler.mreg_14\[24\] _05540_ VGND VGND VPWR VPWR _05541_
+ sky130_fd_sc_hd__xnor2_2
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ clknet_leaf_105_clk _01015_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12693_ _06326_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__clkbuf_1
X_11644_ _05473_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__xor2_2
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ clknet_leaf_96_clk _00946_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput27 hash[123] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
XFILLER_128_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 hash[113] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_14363_ clknet_leaf_15_clk _00877_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11575_ _04762_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__nor2_1
Xinput38 hash[133] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_4
X_10526_ sha256cu.msg_scheduler.mreg_8\[4\] _04526_ _04536_ _04530_ VGND VGND VPWR
+ VPWR _00720_ sky130_fd_sc_hd__o211a_1
X_14294_ clknet_leaf_25_clk _00840_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 hash[143] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
X_13314_ _06656_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10457_ sha256cu.msg_scheduler.mreg_8\[7\] _04494_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__or2_1
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13245_ _06620_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10388_ sha256cu.msg_scheduler.mreg_7\[9\] _04455_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__or2_1
XFILLER_97_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13176_ _06583_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12127_ _05934_ _05937_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12058_ sha256cu.msg_scheduler.mreg_1\[27\] _05870_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11009_ sha256cu.m_pad_pars.m_size\[4\] sha256cu.m_pad_pars.block_512\[63\]\[4\]
+ _01919_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__mux2_1
XFILLER_93_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_290 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08220_ _02824_ _02826_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__and2_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08151_ _02758_ _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__xnor2_2
XFILLER_146_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08082_ sha256cu.K\[17\] _02657_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__a21bo_1
X_07102_ _01622_ _01647_ _01710_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__a21oi_1
X_07033_ _01682_ _01706_ _01652_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08984_ _03472_ _03473_ _03474_ _03366_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__o211a_1
XFILLER_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07935_ sha256cu.m_out_digest.a_in\[14\] _02037_ _02017_ _02550_ VGND VGND VPWR VPWR
+ _02551_ sky130_fd_sc_hd__a22o_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07866_ sha256cu.K\[12\] _02466_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__nand2_1
X_09605_ sha256cu.m_out_digest.g_in\[9\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[9\]
+ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__a22o_1
XFILLER_84_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06817_ net161 net164 net163 net166 VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__or4_1
X_07797_ sha256cu.m_out_digest.e_in\[17\] sha256cu.m_out_digest.e_in\[4\] VGND VGND
+ VPWR VPWR _02416_ sky130_fd_sc_hd__xnor2_2
XFILLER_83_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09536_ _03954_ _03984_ _03980_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__a21o_1
X_09467_ _03936_ _03940_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__nor2_1
X_08418_ _02977_ _02979_ _03020_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__o21ba_1
XFILLER_24_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09398_ _02931_ _03843_ _03844_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__a21boi_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08349_ _02888_ _02916_ _02914_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__o21a_1
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11360_ sha256cu.m_pad_pars.block_512\[5\]\[4\] _05160_ _05161_ sha256cu.m_pad_pars.block_512\[53\]\[4\]
+ _05206_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__a221o_1
XFILLER_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10311_ sha256cu.msg_scheduler.mreg_5\[8\] _04407_ _04413_ _04410_ VGND VGND VPWR
+ VPWR _00628_ sky130_fd_sc_hd__o211a_1
XFILLER_138_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13030_ _06505_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__clkbuf_1
X_11291_ sha256cu.m_pad_pars.block_512\[25\]\[0\] _05140_ _05141_ sha256cu.m_pad_pars.block_512\[29\]\[0\]
+ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__a22o_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10242_ _04281_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__clkbuf_2
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10173_ _04281_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__clkbuf_2
XFILLER_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13932_ clknet_leaf_52_clk _00478_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13863_ clknet_leaf_22_clk _00409_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13794_ clknet_leaf_85_clk _00340_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_12814_ sha256cu.m_pad_pars.block_512\[27\]\[1\] _06389_ VGND VGND VPWR VPWR _06391_
+ sky130_fd_sc_hd__and2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _06354_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _06317_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11627_ _05456_ _05458_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__xnor2_1
X_14415_ clknet_leaf_15_clk _00929_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14346_ clknet_leaf_112_clk _00860_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11558_ sha256cu.m_pad_pars.block_512\[32\]\[7\] _05393_ _04909_ VGND VGND VPWR VPWR
+ _05394_ sky130_fd_sc_hd__o21a_1
XFILLER_144_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10509_ _04447_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__buf_2
X_14277_ clknet_leaf_27_clk _00823_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11489_ sha256cu.m_pad_pars.block_512\[4\]\[1\] _05313_ _05288_ sha256cu.m_pad_pars.block_512\[48\]\[1\]
+ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__a22o_1
XFILLER_143_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13228_ _06611_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13159_ _06574_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__clkbuf_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _02339_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__and2b_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07651_ _02273_ sha256cu.m_out_digest.a_in\[9\] VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__xnor2_4
XFILLER_26_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07582_ _02166_ _02168_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__nor2_1
XFILLER_81_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09321_ _03793_ _03798_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__and2_1
XFILLER_34_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09252_ _02747_ _03696_ _03697_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__a21boi_1
X_09183_ _03664_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__xnor2_1
X_08203_ sha256cu.m_out_digest.e_in\[28\] _02810_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__xnor2_4
XFILLER_147_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08134_ _02026_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__xnor2_2
XFILLER_147_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08065_ _02273_ sha256cu.m_out_digest.a_in\[8\] VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07016_ _01625_ _01643_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__nand2_2
XFILLER_102_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput217 hash[64] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput206 hash[54] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_4
Xinput239 hash[84] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_2
XFILLER_130_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08967_ sha256cu.iter_processing.w\[11\] _02413_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__or2_1
XFILLER_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput228 hash[74] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_2
X_08898_ _03389_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__xnor2_1
X_07918_ _02523_ _02533_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__xor2_1
X_07849_ sha256cu.K\[12\] _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10860_ sha256cu.m_pad_pars.add_out3\[4\] _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__or2_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09519_ _03988_ _03989_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__nand2_1
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10791_ sha256cu.msg_scheduler.mreg_12\[23\] _04679_ VGND VGND VPWR VPWR _04687_
+ sky130_fd_sc_hd__or2_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _06238_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12461_ sha256cu.m_pad_pars.block_512\[6\]\[5\] _06196_ VGND VGND VPWR VPWR _06202_
+ sky130_fd_sc_hd__and2_1
X_14200_ clknet_leaf_28_clk _00746_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_11412_ _04698_ _04801_ _04973_ _05255_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__a31o_1
XFILLER_153_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14131_ clknet_leaf_33_clk _00677_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_12392_ _06165_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11343_ sha256cu.m_pad_pars.block_512\[13\]\[3\] _05128_ _05144_ sha256cu.m_pad_pars.block_512\[9\]\[3\]
+ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__a22o_1
XFILLER_153_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14062_ clknet_leaf_38_clk _00608_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11274_ sha256cu.m_pad_pars.add_out1\[4\] sha256cu.m_pad_pars.add_out1\[5\] VGND
+ VGND VPWR VPWR _05125_ sky130_fd_sc_hd__nor2b_2
X_10225_ sha256cu.msg_scheduler.mreg_4\[3\] _04354_ _04364_ _04357_ VGND VGND VPWR
+ VPWR _00591_ sky130_fd_sc_hd__o211a_1
X_13013_ _06496_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__clkbuf_1
X_10156_ sha256cu.msg_scheduler.mreg_3\[5\] _04315_ _04325_ _04318_ VGND VGND VPWR
+ VPWR _00561_ sky130_fd_sc_hd__o211a_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10087_ sha256cu.msg_scheduler.mreg_3\[8\] _04282_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__or2_1
XFILLER_48_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13915_ clknet_leaf_45_clk _00461_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14895_ clknet_leaf_0_clk _01409_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[59\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13846_ clknet_leaf_17_clk _00392_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13777_ clknet_leaf_66_clk _00323_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10989_ sha256cu.m_pad_pars.block_512\[59\]\[2\] _04829_ VGND VGND VPWR VPWR _04854_
+ sky130_fd_sc_hd__and2_1
X_12728_ sha256cu.m_pad_pars.block_512\[22\]\[1\] _06343_ VGND VGND VPWR VPWR _06345_
+ sky130_fd_sc_hd__and2_1
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12659_ _06308_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14329_ clknet_leaf_90_clk _00024_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09870_ sha256cu.msg_scheduler.mreg_12\[20\] _04153_ _04159_ _04157_ VGND VGND VPWR
+ VPWR _00435_ sky130_fd_sc_hd__o211a_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03296_ _03300_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__nor2_1
XFILLER_112_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _03244_ _03250_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__xor2_1
XFILLER_100_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07703_ _02252_ _02290_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__nor2_1
X_08683_ sha256cu.m_out_digest.d_in\[25\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[25\]
+ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__a22o_1
XFILLER_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07634_ _02002_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__buf_4
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07565_ sha256cu.m_out_digest.g_in\[5\] sha256cu.m_out_digest.f_in\[5\] sha256cu.m_out_digest.e_in\[5\]
+ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__mux2_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07496_ _02121_ _02122_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__and2b_1
X_09304_ _03781_ _03782_ _03779_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09235_ _03715_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__nand2_1
XFILLER_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09166_ sha256cu.iter_processing.w\[18\] _02671_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__nor2_1
XFILLER_134_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09097_ _03582_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__or2_1
X_08117_ _02702_ _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__xor2_1
XFILLER_135_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08048_ _02659_ _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__or2_2
XFILLER_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10010_ sha256cu.msg_scheduler.mreg_2\[7\] _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__or2_1
XFILLER_115_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09999_ sha256cu.msg_scheduler.mreg_1\[2\] _04234_ _04235_ _04224_ VGND VGND VPWR
+ VPWR _00494_ sky130_fd_sc_hd__o211a_1
XFILLER_89_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11961_ _05776_ _05777_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__nand2_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13700_ clknet_leaf_85_clk _00246_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[23\]
+ sky130_fd_sc_hd__dfxtp_4
X_10912_ _04752_ _04776_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__or2_2
X_11892_ sha256cu.msg_scheduler.mreg_9\[13\] sha256cu.msg_scheduler.mreg_0\[13\] VGND
+ VGND VPWR VPWR _05712_ sky130_fd_sc_hd__nand2_1
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14680_ clknet_leaf_119_clk _01194_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[32\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13631_ clknet_leaf_84_clk _00177_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10843_ sha256cu.m_pad_pars.add_out2\[3\] sha256cu.m_pad_pars.add_out2\[2\] VGND
+ VGND VPWR VPWR _04720_ sky130_fd_sc_hd__nand2_1
XFILLER_13_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13562_ clknet_leaf_64_clk _00108_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10774_ sha256cu.msg_scheduler.mreg_11\[15\] _04672_ _04677_ _04675_ VGND VGND VPWR
+ VPWR _00827_ sky130_fd_sc_hd__o211a_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12513_ _06229_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13493_ sha256cu.counter_iteration\[6\] _00051_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__and2b_1
XFILLER_138_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12444_ sha256cu.m_pad_pars.block_512\[5\]\[5\] _06187_ VGND VGND VPWR VPWR _06193_
+ sky130_fd_sc_hd__and2_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12375_ sha256cu.m_pad_pars.block_512\[1\]\[4\] _06152_ VGND VGND VPWR VPWR _06157_
+ sky130_fd_sc_hd__and2_1
X_14114_ clknet_leaf_37_clk _00660_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11326_ sha256cu.m_pad_pars.block_512\[53\]\[1\] _05161_ _05175_ _05024_ VGND VGND
+ VPWR VPWR _05176_ sky130_fd_sc_hd__a22o_1
X_14045_ clknet_leaf_41_clk _00591_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11257_ _01952_ _05004_ _05005_ sha256cu.m_pad_pars.block_512\[50\]\[7\] VGND VGND
+ VPWR VPWR _05109_ sky130_fd_sc_hd__o22a_1
X_10208_ sha256cu.msg_scheduler.mreg_4\[28\] _04348_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__or2_1
XFILLER_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11188_ sha256cu.m_pad_pars.block_512\[6\]\[3\] _04957_ _04989_ sha256cu.m_pad_pars.block_512\[14\]\[3\]
+ _05043_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__a221o_1
X_10139_ sha256cu.msg_scheduler.mreg_3\[30\] _04308_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__or2_1
XFILLER_79_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14947_ clknet_leaf_91_clk _01461_ VGND VGND VPWR VPWR sha256cu.K\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_62_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14878_ clknet_leaf_117_clk _01392_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13829_ clknet_leaf_109_clk _00375_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[24\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_62_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07350_ sha256cu.m_pad_pars.add_out0\[2\] _01963_ _01966_ VGND VGND VPWR VPWR _01990_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09020_ _03507_ _03508_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__nor2_1
XFILLER_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07281_ sha256cu.m_pad_pars.m_size\[4\] sha256cu.m_pad_pars.block_512\[63\]\[4\]
+ _01928_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__mux2_1
XFILLER_129_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09922_ sha256cu.msg_scheduler.mreg_1\[1\] _04174_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__or2_1
XFILLER_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09853_ sha256cu.msg_scheduler.mreg_13\[13\] _04147_ VGND VGND VPWR VPWR _04150_
+ sky130_fd_sc_hd__or2_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _03296_ _03300_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__xor2_1
XFILLER_112_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09784_ sha256cu.msg_scheduler.mreg_14\[16\] _04106_ VGND VGND VPWR VPWR _04110_
+ sky130_fd_sc_hd__or2_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _03232_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__xor2_1
XFILLER_65_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _01590_ _01633_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__nor2_4
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ sha256cu.m_out_digest.d_in\[10\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[10\]
+ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__o22a_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07617_ _02228_ _02240_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__xor2_2
XFILLER_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ sha256cu.m_out_digest.b_in\[17\] _03177_ _03176_ _02162_ VGND VGND VPWR VPWR
+ _00144_ sky130_fd_sc_hd__o22a_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07548_ _02150_ _02173_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07479_ sha256cu.m_out_digest.a_in\[2\] _02002_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__or2_1
XFILLER_50_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10490_ _04396_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__buf_2
X_09218_ _02712_ _03671_ _03672_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a21boi_1
XFILLER_10_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09149_ _03632_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12160_ sha256cu.msg_scheduler.mreg_9\[24\] sha256cu.msg_scheduler.mreg_0\[24\] VGND
+ VGND VPWR VPWR _05969_ sky130_fd_sc_hd__nand2_1
Xpassword_cracker_262 VGND VGND VPWR VPWR password_cracker_262/HI password_count[2]
+ sky130_fd_sc_hd__conb_1
Xpassword_cracker_284 VGND VGND VPWR VPWR password_cracker_284/HI password_count[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11111_ _04797_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__inv_2
XFILLER_2_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpassword_cracker_273 VGND VGND VPWR VPWR password_cracker_273/HI password_count[13]
+ sky130_fd_sc_hd__conb_1
X_12091_ _05900_ _05901_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__and2_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11042_ _04897_ _04898_ _04900_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__or4_2
XFILLER_103_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14801_ clknet_leaf_1_clk _01315_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12993_ sha256cu.m_pad_pars.block_512\[37\]\[5\] _06480_ VGND VGND VPWR VPWR _06486_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11944_ _05760_ _05761_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__nor2_1
X_14732_ clknet_leaf_7_clk _01246_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11875_ _05693_ _05694_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__nand2_1
X_14663_ clknet_leaf_13_clk _01177_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[30\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13614_ clknet_leaf_73_clk _00160_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10826_ sha256cu.m_pad_pars.add_512_block\[2\] _04700_ _04710_ _04709_ VGND VGND
+ VPWR VPWR _00846_ sky130_fd_sc_hd__o211a_1
XFILLER_60_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14594_ clknet_leaf_101_clk _01108_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10757_ sha256cu.msg_scheduler.mreg_12\[8\] _04666_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__or2_1
X_13545_ clknet_leaf_79_clk _00091_ VGND VGND VPWR VPWR Hash_Digest sky130_fd_sc_hd__dfxtp_1
XFILLER_41_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10688_ sha256cu.msg_scheduler.mreg_11\[10\] _04627_ VGND VGND VPWR VPWR _04629_
+ sky130_fd_sc_hd__or2_1
X_13476_ _06749_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12427_ sha256cu.m_pad_pars.block_512\[4\]\[5\] _06178_ VGND VGND VPWR VPWR _06184_
+ sky130_fd_sc_hd__and2_1
XFILLER_126_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12358_ _06148_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12289_ _06072_ _06075_ _06092_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__o21ai_1
X_11309_ _04768_ _05159_ _05152_ _05127_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__o211a_2
X_14028_ clknet_leaf_56_clk _00574_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06850_ _01544_ _01545_ _01546_ _01547_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__or4_1
XFILLER_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06781_ net78 net111 net100 net134 VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__or4_4
X_08520_ _03117_ _03119_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__xnor2_1
X_08451_ _03051_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__xnor2_1
X_07402_ _02022_ _02031_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__nor2_1
XFILLER_63_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08382_ _02984_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__or2_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07333_ _01964_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_124_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_32_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07264_ sha256cu.byte_rdy sha256cu.byte_stop VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__or2b_1
X_09003_ _03491_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__xor2_1
XFILLER_3_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07195_ _01647_ _01610_ _01706_ _01859_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__a31o_1
XFILLER_145_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09905_ sha256cu.msg_scheduler.counter_iteration\[3\] sha256cu.msg_scheduler.counter_iteration\[2\]
+ _04178_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__and3_1
XFILLER_101_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09836_ _04044_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__buf_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09767_ sha256cu.msg_scheduler.mreg_13\[8\] _04099_ _04100_ _04090_ VGND VGND VPWR
+ VPWR _00391_ sky130_fd_sc_hd__o211a_1
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06979_ _01577_ _00453_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__nor2_4
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _03193_ _03196_ _03217_ _02923_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__a31oi_1
X_09698_ sha256cu.msg_scheduler.mreg_14\[10\] _04060_ _04061_ _04050_ VGND VGND VPWR
+ VPWR _00361_ sky130_fd_sc_hd__o211a_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ sha256cu.m_out_digest.c_in\[29\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[29\]
+ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__o22a_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11660_ _05487_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__xor2_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ sha256cu.msg_scheduler.mreg_9\[8\] _04581_ _04585_ _04584_ VGND VGND VPWR
+ VPWR _00756_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_115_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_16
X_11591_ _05398_ _05403_ _05409_ _05426_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__or4_1
X_10542_ sha256cu.msg_scheduler.mreg_8\[11\] _04540_ _04545_ _04543_ VGND VGND VPWR
+ VPWR _00727_ sky130_fd_sc_hd__o211a_1
X_13330_ sha256cu.m_pad_pars.block_512\[57\]\[3\] _06660_ VGND VGND VPWR VPWR _06665_
+ sky130_fd_sc_hd__and2_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13261_ sha256cu.m_pad_pars.block_512\[53\]\[2\] _06626_ VGND VGND VPWR VPWR _06629_
+ sky130_fd_sc_hd__and2_1
XFILLER_10_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10473_ sha256cu.msg_scheduler.mreg_8\[14\] _04494_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__or2_1
X_12212_ _06017_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__and2_1
XFILLER_41_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13192_ _06592_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_1
X_12143_ _05923_ _05927_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__nand3_1
XFILLER_151_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12074_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__inv_2
XFILLER_150_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11025_ sha256cu.m_pad_pars.block_512\[27\]\[5\] _04757_ _04804_ sha256cu.m_pad_pars.block_512\[43\]\[5\]
+ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__a221o_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14715_ clknet_leaf_125_clk _01229_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12976_ sha256cu.m_pad_pars.block_512\[36\]\[5\] _06471_ VGND VGND VPWR VPWR _06477_
+ sky130_fd_sc_hd__and2_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _05720_ _05722_ _05718_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__a21oi_1
XFILLER_72_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _05677_ _05679_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14646_ clknet_leaf_113_clk _01160_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10809_ sha256cu.msg_scheduler.mreg_12\[31\] _04692_ VGND VGND VPWR VPWR _04697_
+ sky130_fd_sc_hd__or2_1
X_11789_ _05612_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__xor2_1
XANTENNA_19 _01994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_106_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_13_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14577_ clknet_leaf_4_clk _01091_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13528_ clknet_leaf_2_clk _00078_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13459_ _04188_ _00037_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__and2b_1
XFILLER_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07951_ _02565_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__inv_2
XFILLER_101_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06902_ _01593_ _01590_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__and3_2
X_07882_ _02451_ _02454_ _02498_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__o21a_1
XFILLER_68_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06833_ net107 net110 net109 net114 VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__or4_1
X_09621_ _02923_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__buf_4
XFILLER_56_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09552_ _04004_ _04007_ _04022_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__and3_1
XFILLER_55_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08503_ _03075_ _03103_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__xnor2_1
X_09483_ sha256cu.m_out_digest.e_in\[28\] _02732_ _03954_ _03956_ _01913_ VGND VGND
+ VPWR VPWR _00251_ sky130_fd_sc_hd__a221o_1
XFILLER_51_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08434_ _02996_ _03022_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__nor2_1
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08365_ sha256cu.m_out_digest.b_in\[26\] _02161_ sha256cu.m_out_digest.c_in\[26\]
+ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__a21o_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07316_ _01949_ _01955_ _01959_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__a21o_1
XFILLER_32_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08296_ sha256cu.m_out_digest.b_in\[24\] _02083_ _02901_ VGND VGND VPWR VPWR _02902_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_07247_ _01752_ _01904_ _01629_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__o21a_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07178_ _01591_ _01612_ _01776_ _01652_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__a211o_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09819_ sha256cu.msg_scheduler.mreg_13\[30\] _04126_ _04129_ _04130_ VGND VGND VPWR
+ VPWR _00413_ sky130_fd_sc_hd__o211a_1
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12830_ _06399_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__clkbuf_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12761_ sha256cu.m_pad_pars.block_512\[24\]\[0\] _06362_ VGND VGND VPWR VPWR _06363_
+ sky130_fd_sc_hd__and2_1
XFILLER_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ sha256cu.msg_scheduler.mreg_14\[22\] sha256cu.msg_scheduler.mreg_14\[15\]
+ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__xnor2_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ sha256cu.m_pad_pars.block_512\[20\]\[0\] _06325_ VGND VGND VPWR VPWR _06326_
+ sky130_fd_sc_hd__and2_1
X_14500_ clknet_leaf_103_clk _01014_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11643_ _05450_ _05453_ _05449_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a21boi_2
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ clknet_leaf_97_clk _00945_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 hash[114] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14362_ clknet_leaf_14_clk _00876_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput28 hash[124] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlymetal6s2s_1
X_11574_ _04786_ _05291_ sha256cu.m_pad_pars.block_512\[4\]\[7\] VGND VGND VPWR VPWR
+ _05410_ sky130_fd_sc_hd__a21oi_1
X_10525_ sha256cu.msg_scheduler.mreg_9\[4\] _04534_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__or2_1
Xinput39 hash[134] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
X_14293_ clknet_leaf_27_clk _00839_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_13313_ sha256cu.m_pad_pars.block_512\[56\]\[3\] _01924_ VGND VGND VPWR VPWR _06656_
+ sky130_fd_sc_hd__and2_1
X_10456_ sha256cu.msg_scheduler.mreg_7\[6\] _04487_ _04496_ _04490_ VGND VGND VPWR
+ VPWR _00690_ sky130_fd_sc_hd__o211a_1
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13244_ sha256cu.m_pad_pars.block_512\[52\]\[2\] _06617_ VGND VGND VPWR VPWR _06620_
+ sky130_fd_sc_hd__and2_1
X_13175_ sha256cu.m_pad_pars.block_512\[48\]\[2\] _06580_ VGND VGND VPWR VPWR _06583_
+ sky130_fd_sc_hd__and2_1
X_10387_ sha256cu.msg_scheduler.mreg_6\[8\] _04448_ _04457_ _04451_ VGND VGND VPWR
+ VPWR _00660_ sky130_fd_sc_hd__o211a_1
X_12126_ _05890_ _05935_ _05936_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__a21bo_1
XFILLER_151_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12057_ sha256cu.msg_scheduler.mreg_1\[23\] sha256cu.msg_scheduler.mreg_1\[6\] VGND
+ VGND VPWR VPWR _05870_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11008_ _01971_ _04870_ _04871_ _04709_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__o211a_1
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12959_ sha256cu.m_pad_pars.block_512\[35\]\[5\] _06462_ VGND VGND VPWR VPWR _06468_
+ sky130_fd_sc_hd__and2_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_291 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_280 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14629_ clknet_leaf_97_clk _01143_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08150_ sha256cu.K\[19\] _02726_ _02759_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__a21oi_2
XFILLER_119_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07101_ _01679_ _01774_ _01778_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__a21o_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08081_ _02656_ _02634_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__or2b_1
X_07032_ _01666_ _01714_ _01715_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08983_ sha256cu.m_out_digest.e_in\[11\] _02440_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__or2_1
X_07934_ _02545_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07865_ _02463_ _02465_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__or2b_1
XFILLER_69_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09604_ sha256cu.m_out_digest.g_in\[8\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[8\]
+ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__o22a_1
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07796_ sha256cu.iter_processing.w\[11\] _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__xnor2_2
X_06816_ net157 net160 net159 net162 VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__or4_2
X_09535_ _03954_ _03984_ _04006_ _03980_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__a211o_1
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09466_ sha256cu.K\[28\] _03939_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__xnor2_1
X_08417_ _02974_ _02976_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__and2b_1
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09397_ _02964_ _03872_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__xor2_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08348_ _02951_ _02952_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__or2_1
X_08279_ _02879_ _02884_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__and2_1
XFILLER_153_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10310_ sha256cu.msg_scheduler.mreg_6\[8\] _04401_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__or2_1
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11290_ _04747_ _05124_ _01977_ _01985_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__o211a_2
XFILLER_153_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10241_ sha256cu.msg_scheduler.mreg_4\[10\] _04367_ _04373_ _04370_ VGND VGND VPWR
+ VPWR _00598_ sky130_fd_sc_hd__o211a_1
XFILLER_98_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10172_ sha256cu.msg_scheduler.mreg_3\[12\] _04328_ _04334_ _04331_ VGND VGND VPWR
+ VPWR _00568_ sky130_fd_sc_hd__o211a_1
XFILLER_79_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13931_ clknet_leaf_52_clk _00477_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13862_ clknet_leaf_23_clk _00408_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13793_ clknet_leaf_84_clk _00339_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[20\]
+ sky130_fd_sc_hd__dfxtp_2
X_12813_ _06390_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12744_ sha256cu.m_pad_pars.block_512\[23\]\[0\] _06353_ VGND VGND VPWR VPWR _06354_
+ sky130_fd_sc_hd__and2_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12675_ sha256cu.m_pad_pars.block_512\[19\]\[0\] _06316_ VGND VGND VPWR VPWR _06317_
+ sky130_fd_sc_hd__and2_1
X_11626_ sha256cu.msg_scheduler.mreg_14\[20\] _05457_ VGND VGND VPWR VPWR _05458_
+ sky130_fd_sc_hd__xnor2_1
X_14414_ clknet_leaf_110_clk _00928_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[30\]
+ sky130_fd_sc_hd__dfxtp_2
X_14345_ clknet_leaf_111_clk _00859_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out3\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_11557_ _04792_ _05136_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__nor2_1
X_10508_ sha256cu.msg_scheduler.mreg_7\[29\] _04513_ _04525_ _04516_ VGND VGND VPWR
+ VPWR _00713_ sky130_fd_sc_hd__o211a_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14276_ clknet_leaf_20_clk _00822_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11488_ sha256cu.m_pad_pars.block_512\[32\]\[1\] _05306_ _05310_ sha256cu.m_pad_pars.block_512\[52\]\[1\]
+ _05329_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__a221o_1
X_10439_ sha256cu.msg_scheduler.mreg_6\[31\] _04474_ _04486_ _04477_ VGND VGND VPWR
+ VPWR _00683_ sky130_fd_sc_hd__o211a_1
X_13227_ sha256cu.m_pad_pars.block_512\[51\]\[2\] _06608_ VGND VGND VPWR VPWR _06611_
+ sky130_fd_sc_hd__and2_1
XFILLER_112_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13158_ sha256cu.m_pad_pars.block_512\[47\]\[2\] _06571_ VGND VGND VPWR VPWR _06574_
+ sky130_fd_sc_hd__and2_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ sha256cu.msg_scheduler.mreg_1\[29\] _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13089_ sha256cu.m_pad_pars.block_512\[43\]\[2\] _06534_ VGND VGND VPWR VPWR _06537_
+ sky130_fd_sc_hd__and2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07650_ sha256cu.m_out_digest.a_in\[20\] VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__buf_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07581_ _02194_ _02205_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__xor2_1
XFILLER_93_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09320_ _03793_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nor2_1
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09251_ _02777_ _03731_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__xor2_1
X_08202_ sha256cu.m_out_digest.e_in\[15\] sha256cu.m_out_digest.e_in\[1\] VGND VGND
+ VPWR VPWR _02810_ sky130_fd_sc_hd__xnor2_4
X_09182_ _03608_ _03638_ _03637_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__a31o_1
X_08133_ sha256cu.m_out_digest.a_in\[10\] sha256cu.m_out_digest.a_in\[1\] VGND VGND
+ VPWR VPWR _02743_ sky130_fd_sc_hd__xnor2_2
XFILLER_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08064_ _02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__inv_2
X_07015_ _01646_ _01680_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__nor2_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput207 hash[55] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput218 hash[65] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_1
Xinput229 hash[75] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_4
X_08966_ _03455_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08897_ _03315_ _03338_ _03362_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__o31a_2
X_07917_ _02530_ _02532_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_95_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
X_07848_ _02463_ _02465_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07779_ _02357_ _02359_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__nor2_1
X_09518_ _03988_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__or2_1
XFILLER_72_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10790_ sha256cu.msg_scheduler.mreg_11\[22\] _04685_ _04686_ _04675_ VGND VGND VPWR
+ VPWR _00834_ sky130_fd_sc_hd__o211a_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ sha256cu.m_out_digest.e_in\[27\] _02439_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__or2_1
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12460_ _06201_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12391_ sha256cu.m_pad_pars.block_512\[2\]\[4\] _06160_ VGND VGND VPWR VPWR _06165_
+ sky130_fd_sc_hd__and2_1
X_11411_ _04917_ _05248_ sha256cu.m_pad_pars.block_512\[45\]\[7\] VGND VGND VPWR VPWR
+ _05255_ sky130_fd_sc_hd__o21a_1
X_14130_ clknet_leaf_34_clk _00676_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11342_ sha256cu.data_in_padd\[18\] _04741_ _04742_ _05190_ VGND VGND VPWR VPWR _00881_
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14061_ clknet_leaf_38_clk _00607_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11273_ _04702_ _01939_ _04776_ sha256cu.m_pad_pars.add_512_block\[1\] VGND VGND
+ VPWR VPWR _05124_ sky130_fd_sc_hd__a211o_2
XFILLER_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10224_ sha256cu.msg_scheduler.mreg_5\[3\] _04361_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__or2_1
X_13012_ sha256cu.m_pad_pars.block_512\[38\]\[6\] _06489_ VGND VGND VPWR VPWR _06496_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10155_ sha256cu.msg_scheduler.mreg_4\[5\] _04322_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__or2_1
XFILLER_133_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10086_ sha256cu.msg_scheduler.mreg_2\[7\] _04274_ _04285_ _04277_ VGND VGND VPWR
+ VPWR _00531_ sky130_fd_sc_hd__o211a_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_48_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13914_ clknet_leaf_46_clk _00460_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14894_ clknet_leaf_9_clk _01408_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13845_ clknet_leaf_17_clk _00391_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13776_ clknet_leaf_66_clk _00322_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10988_ sha256cu.m_pad_pars.block_512\[31\]\[2\] _04811_ _04822_ sha256cu.m_pad_pars.block_512\[47\]\[2\]
+ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__a22o_1
XFILLER_95_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12727_ _06344_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12658_ sha256cu.m_pad_pars.block_512\[18\]\[0\] _06307_ VGND VGND VPWR VPWR _06308_
+ sky130_fd_sc_hd__and2_1
XFILLER_129_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11609_ sha256cu.flag_0_15 sha256cu.msg_scheduler.counter_iteration\[6\] sha256cu.msg_scheduler.counter_iteration\[5\]
+ _05431_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__or4_4
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12589_ _06270_ _04988_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_10_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14328_ clknet_leaf_90_clk _00023_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14259_ clknet_leaf_26_clk _00805_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03294_ _03295_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__nor2_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _03248_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_77_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07702_ _02104_ _02146_ _02181_ _02215_ _02145_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__o2111a_1
X_08682_ sha256cu.m_out_digest.d_in\[24\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[24\]
+ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__o22a_1
X_07633_ _02252_ _02255_ _02069_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07564_ sha256cu.m_out_digest.b_in\[5\] sha256cu.m_out_digest.a_in\[5\] sha256cu.m_out_digest.c_in\[5\]
+ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__a21o_1
XFILLER_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07495_ _02118_ _02119_ _02120_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__a21o_1
X_09303_ _03779_ _03781_ _03782_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__or3_1
X_09234_ _03686_ _03687_ _03684_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__a21o_1
X_09165_ _03647_ _03648_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08116_ sha256cu.K\[19\] _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__xnor2_2
XFILLER_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09096_ _03551_ _03557_ _03581_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__a21oi_1
X_08047_ _02632_ _02617_ _02658_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__a21oi_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09998_ sha256cu.msg_scheduler.mreg_2\[2\] _04228_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__or2_1
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08949_ _03421_ _03422_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__a21o_1
XFILLER_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11960_ sha256cu.msg_scheduler.mreg_9\[16\] sha256cu.msg_scheduler.mreg_0\[16\] VGND
+ VGND VPWR VPWR _05777_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_68_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10911_ _04775_ _04777_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__nand2_1
XFILLER_45_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11891_ sha256cu.msg_scheduler.mreg_9\[13\] sha256cu.msg_scheduler.mreg_0\[13\] VGND
+ VGND VPWR VPWR _05711_ sky130_fd_sc_hd__or2_1
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13630_ clknet_leaf_69_clk _00176_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10842_ _04718_ _04719_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__nor2_1
XFILLER_60_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13561_ clknet_leaf_64_clk _00107_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10773_ sha256cu.msg_scheduler.mreg_12\[15\] _04666_ VGND VGND VPWR VPWR _04677_
+ sky130_fd_sc_hd__or2_1
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12512_ sha256cu.m_pad_pars.block_512\[9\]\[5\] _06223_ VGND VGND VPWR VPWR _06229_
+ sky130_fd_sc_hd__and2_1
XFILLER_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13492_ _06759_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12443_ _06192_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12374_ _06156_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14113_ clknet_leaf_37_clk _00659_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11325_ sha256cu.m_pad_pars.block_512\[61\]\[1\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[1\]
+ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__a22o_1
XFILLER_153_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14044_ clknet_leaf_42_clk _00590_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11256_ _04747_ _04993_ _05107_ sha256cu.m_pad_pars.block_512\[18\]\[7\] VGND VGND
+ VPWR VPWR _05108_ sky130_fd_sc_hd__o22a_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10207_ _04314_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__buf_2
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11187_ sha256cu.m_pad_pars.block_512\[2\]\[3\] _04999_ _05042_ _01921_ VGND VGND
+ VPWR VPWR _05043_ sky130_fd_sc_hd__a22o_1
X_10138_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__buf_2
XFILLER_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_59_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
X_10069_ sha256cu.msg_scheduler.mreg_2\[0\] _04274_ _04275_ _04264_ VGND VGND VPWR
+ VPWR _00524_ sky130_fd_sc_hd__o211a_1
XFILLER_85_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14946_ clknet_leaf_91_clk _01460_ VGND VGND VPWR VPWR sha256cu.K\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14877_ clknet_leaf_125_clk _01391_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13828_ clknet_leaf_110_clk _00374_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[23\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13759_ clknet_leaf_69_clk _00305_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07280_ _01929_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09921_ sha256cu.msg_scheduler.mreg_0\[0\] _04167_ _04191_ _04171_ VGND VGND VPWR
+ VPWR _00460_ sky130_fd_sc_hd__o211a_1
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09852_ sha256cu.msg_scheduler.mreg_12\[12\] _04140_ _04149_ _04144_ VGND VGND VPWR
+ VPWR _00427_ sky130_fd_sc_hd__o211a_1
XFILLER_86_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ sha256cu.K\[5\] _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__xor2_1
XFILLER_112_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09783_ sha256cu.msg_scheduler.mreg_13\[15\] _04099_ _04109_ _04103_ VGND VGND VPWR
+ VPWR _00398_ sky130_fd_sc_hd__o211a_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08734_ _03210_ _03215_ _03233_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__o21ai_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _01648_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__and2_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ sha256cu.m_out_digest.d_in\[9\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[9\]
+ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__a22o_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07616_ _02237_ _02239_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__xnor2_2
XFILLER_121_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _02369_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__buf_4
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07547_ _02170_ _02172_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07478_ _02104_ _02105_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__or2_1
XFILLER_10_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09217_ _02747_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__xor2_1
XFILLER_148_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09148_ sha256cu.K\[16\] _03595_ _03594_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__a21o_1
X_09079_ _03564_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__nor2_1
Xpassword_cracker_263 VGND VGND VPWR VPWR password_cracker_263/HI password_count[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_150_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpassword_cracker_274 VGND VGND VPWR VPWR password_cracker_274/HI password_count[14]
+ sky130_fd_sc_hd__conb_1
Xpassword_cracker_285 VGND VGND VPWR VPWR password_cracker_285/HI password_count[25]
+ sky130_fd_sc_hd__conb_1
X_11110_ _04704_ _04954_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__or2_2
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12090_ _05900_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__nor2_1
XFILLER_131_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11041_ sha256cu.m_pad_pars.block_512\[3\]\[6\] _04765_ _04826_ sha256cu.m_pad_pars.block_512\[51\]\[6\]
+ _04901_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__a221o_1
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14800_ clknet_leaf_0_clk _01314_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[47\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12992_ _06485_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11943_ _05731_ _05735_ _05732_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a21boi_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14731_ clknet_leaf_8_clk _01245_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11874_ _05693_ _05694_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__or2_1
XFILLER_72_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14662_ clknet_leaf_116_clk _01176_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13613_ clknet_leaf_74_clk _00159_ VGND VGND VPWR VPWR sha256cu.m_out_digest.c_in\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10825_ sha256cu.m_pad_pars.m_size\[5\] _04706_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__or2_1
X_14593_ clknet_leaf_104_clk _01107_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10756_ sha256cu.msg_scheduler.mreg_11\[7\] _04659_ _04667_ _04662_ VGND VGND VPWR
+ VPWR _00819_ sky130_fd_sc_hd__o211a_1
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13544_ clknet_leaf_105_clk _00090_ VGND VGND VPWR VPWR sha256cu.iter_processing.temp_if
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10687_ sha256cu.msg_scheduler.mreg_10\[9\] _04620_ _04628_ _04623_ VGND VGND VPWR
+ VPWR _00789_ sky130_fd_sc_hd__o211a_1
XFILLER_9_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13475_ _06730_ _06748_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__and2_1
XFILLER_139_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12426_ _06183_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__clkbuf_1
X_12357_ sha256cu.m_pad_pars.block_512\[0\]\[3\] _06144_ VGND VGND VPWR VPWR _06148_
+ sky130_fd_sc_hd__and2_1
XFILLER_141_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12288_ _06090_ _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__and2b_1
X_11308_ sha256cu.m_pad_pars.temp_chk _04954_ _05154_ sha256cu.m_pad_pars.add_512_block\[6\]
+ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__o22a_2
X_14027_ clknet_leaf_56_clk _00573_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11239_ _04768_ _04960_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__or2_1
XFILLER_110_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06780_ net245 net23 net12 net45 VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__or4_2
XFILLER_83_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14929_ clknet_leaf_95_clk _01443_ VGND VGND VPWR VPWR sha256cu.K\[2\] sky130_fd_sc_hd__dfxtp_2
X_08450_ sha256cu.m_out_digest.g_in\[28\] sha256cu.m_out_digest.f_in\[28\] sha256cu.m_out_digest.e_in\[28\]
+ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__mux2_2
X_07401_ _02025_ _02030_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08381_ _02981_ _02982_ sha256cu.K\[26\] VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__and3b_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07332_ sha256cu.m_pad_pars.add_out1\[3\] _01962_ _01968_ _01971_ _01974_ VGND VGND
+ VPWR VPWR _00082_ sky130_fd_sc_hd__o221a_1
XFILLER_149_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07263_ _01914_ _01915_ sha256cu.m_pad_pars.add_512_block\[6\] VGND VGND VPWR VPWR
+ _01916_ sky130_fd_sc_hd__a21oi_2
X_09002_ sha256cu.K\[11\] _03458_ _03459_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__a21bo_1
X_07194_ _01622_ _01603_ _01652_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09904_ sha256cu.msg_scheduler.counter_iteration\[2\] _04178_ _04180_ VGND VGND VPWR
+ VPWR _00448_ sky130_fd_sc_hd__o21a_1
XFILLER_98_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09835_ sha256cu.msg_scheduler.mreg_12\[5\] _04126_ _04139_ _04130_ VGND VGND VPWR
+ VPWR _00420_ sky130_fd_sc_hd__o211a_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09766_ sha256cu.msg_scheduler.mreg_14\[8\] _04093_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__or2_1
XFILLER_86_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06978_ _00454_ _01665_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__nand2_4
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _03193_ _03196_ _03217_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__a21o_1
X_09697_ sha256cu.iter_processing.w\[10\] _04054_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__or2_1
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ sha256cu.m_out_digest.c_in\[28\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[28\]
+ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__o22a_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ sha256cu.m_out_digest.b_in\[1\] _03031_ _02114_ sha256cu.m_out_digest.a_in\[1\]
+ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__a22o_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ sha256cu.msg_scheduler.mreg_10\[8\] _04574_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__or2_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11590_ _05412_ _05418_ _05422_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__or4b_1
XFILLER_128_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10541_ sha256cu.msg_scheduler.mreg_9\[11\] _04534_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__or2_1
X_13260_ _06628_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10472_ sha256cu.msg_scheduler.mreg_7\[13\] _04500_ _04505_ _04503_ VGND VGND VPWR
+ VPWR _00697_ sky130_fd_sc_hd__o211a_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12211_ _06015_ _06016_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__nand2_1
XFILLER_6_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13191_ sha256cu.m_pad_pars.block_512\[49\]\[1\] _06590_ VGND VGND VPWR VPWR _06592_
+ sky130_fd_sc_hd__and2_1
XFILLER_150_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12142_ _05950_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12073_ _05840_ _05819_ _05860_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__nand3b_1
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11024_ sha256cu.m_pad_pars.block_512\[51\]\[5\] _04826_ _04822_ sha256cu.m_pad_pars.block_512\[47\]\[5\]
+ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__a221o_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12975_ _06476_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11926_ _05743_ _05744_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__nand2_1
XFILLER_80_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14714_ clknet_leaf_126_clk _01228_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ sha256cu.msg_scheduler.mreg_14\[30\] _05678_ VGND VGND VPWR VPWR _05679_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_60_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14645_ clknet_leaf_3_clk _01159_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11788_ _05579_ _05581_ _05577_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__a21oi_1
X_10808_ sha256cu.msg_scheduler.mreg_11\[30\] _04685_ _04696_ _04688_ VGND VGND VPWR
+ VPWR _00842_ sky130_fd_sc_hd__o211a_1
X_14576_ clknet_leaf_2_clk _01090_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10739_ sha256cu.msg_scheduler.mreg_11\[0\] _04646_ _04657_ _04649_ VGND VGND VPWR
+ VPWR _00812_ sky130_fd_sc_hd__o211a_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13527_ clknet_leaf_124_clk _00077_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13458_ sha256cu.K\[9\] _06726_ _06727_ _06738_ _06737_ VGND VGND VPWR VPWR _01450_
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12409_ _06174_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__clkbuf_1
X_13389_ sha256cu.m_pad_pars.block_512\[60\]\[7\] _06693_ VGND VGND VPWR VPWR _06696_
+ sky130_fd_sc_hd__and2_1
XFILLER_102_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07950_ sha256cu.m_out_digest.e_in\[26\] _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__xnor2_2
XFILLER_141_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06901_ _01592_ _00452_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__or2_2
X_07881_ sha256cu.m_out_digest.h_in\[12\] _02453_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__nand2_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06832_ net103 net106 net105 net108 VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__or4_1
X_09620_ sha256cu.m_out_digest.g_in\[21\] _04033_ _04036_ sha256cu.m_out_digest.f_in\[21\]
+ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__a22o_1
XFILLER_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09551_ _04015_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08502_ _03101_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__or2b_1
XFILLER_102_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09482_ _02629_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__nor2_1
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08433_ _03019_ _03021_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__nor2_1
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08364_ _02965_ _02967_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07315_ _01919_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__and2_1
XFILLER_149_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08295_ sha256cu.m_out_digest.b_in\[24\] _02083_ sha256cu.m_out_digest.c_in\[24\]
+ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__a21o_1
X_07246_ _01613_ _01695_ _01644_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07177_ _01621_ _01844_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__or2_1
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09818_ _04116_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__buf_2
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09749_ sha256cu.msg_scheduler.mreg_13\[0\] _04086_ _04089_ _04090_ VGND VGND VPWR
+ VPWR _00383_ sky130_fd_sc_hd__o211a_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _06251_ _05081_ _05276_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__or3_4
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _05537_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__and2b_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _06251_ _05081_ _05292_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__or3_4
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11642_ _05470_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__xor2_2
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14430_ clknet_leaf_116_clk _00944_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14361_ clknet_leaf_14_clk _00875_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 hash[115] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
XFILLER_11_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13312_ _06655_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
X_11573_ _05278_ _05277_ _05405_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__a31o_1
X_10524_ sha256cu.msg_scheduler.mreg_8\[3\] _04526_ _04535_ _04530_ VGND VGND VPWR
+ VPWR _00719_ sky130_fd_sc_hd__o211a_1
Xinput29 hash[125] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
X_14292_ clknet_leaf_25_clk _00838_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10455_ sha256cu.msg_scheduler.mreg_8\[6\] _04494_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__or2_1
XFILLER_109_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13243_ _06619_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13174_ _06582_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10386_ sha256cu.msg_scheduler.mreg_7\[8\] _04455_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__or2_1
X_12125_ _05883_ _05909_ _05908_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__a21o_1
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12056_ _05867_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nand2_1
XFILLER_93_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11007_ sha256cu.data_in_padd\[3\] _01963_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__or2_1
XFILLER_92_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12958_ _06467_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ _05727_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__nor2_1
XFILLER_61_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12889_ _06430_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_270 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_292 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14628_ clknet_leaf_97_clk _01142_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_281 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07100_ _01595_ _01729_ _01775_ _01777_ _01629_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__o311a_1
X_14559_ clknet_leaf_96_clk _01073_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_08080_ sha256cu.K\[18\] _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__xnor2_2
X_07031_ _01643_ _01639_ _01680_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__and3_1
XFILLER_130_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08982_ _03441_ _03448_ _03471_ _02629_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a31o_1
X_07933_ _02476_ _02547_ _02548_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__o21bai_1
XFILLER_69_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07864_ _02467_ _02469_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__and2b_1
XFILLER_69_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09603_ sha256cu.m_out_digest.g_in\[7\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[7\]
+ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__o22a_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06815_ net148 net151 net150 net153 VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__or4_2
X_07795_ _02412_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__xnor2_2
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09534_ _04004_ _04005_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__nand2_1
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09465_ _03937_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__nor2_1
XFILLER_36_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08416_ _03016_ _03018_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09396_ _03870_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__nand2_1
X_08347_ _02924_ _02950_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__nor2_1
XFILLER_138_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08278_ _02766_ _02878_ _02880_ _02883_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__o211a_1
XFILLER_20_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07229_ _01632_ _01615_ _01673_ _01618_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__o211a_1
X_10240_ sha256cu.msg_scheduler.mreg_5\[10\] _04361_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__or2_1
XFILLER_106_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10171_ sha256cu.msg_scheduler.mreg_4\[12\] _04322_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__or2_1
XFILLER_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13930_ clknet_leaf_52_clk _00476_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13861_ clknet_leaf_23_clk _00407_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13792_ clknet_leaf_84_clk _00338_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12812_ sha256cu.m_pad_pars.block_512\[27\]\[0\] _06389_ VGND VGND VPWR VPWR _06390_
+ sky130_fd_sc_hd__and2_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12743_ _01912_ _04827_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__or2_2
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ clknet_leaf_110_clk _00927_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[29\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _01912_ _04830_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__or2_2
XFILLER_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11625_ sha256cu.msg_scheduler.mreg_14\[18\] sha256cu.msg_scheduler.mreg_14\[11\]
+ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14344_ clknet_leaf_112_clk _00858_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out3\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_7_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11556_ _01992_ _05391_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__and2_1
X_10507_ sha256cu.msg_scheduler.mreg_8\[29\] _04520_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__or2_1
X_14275_ clknet_leaf_20_clk _00821_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13226_ _06610_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
X_11487_ sha256cu.m_pad_pars.block_512\[44\]\[1\] _05298_ _05296_ sha256cu.m_pad_pars.block_512\[28\]\[1\]
+ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__a22o_1
X_10438_ sha256cu.msg_scheduler.mreg_7\[31\] _04481_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__or2_1
XFILLER_152_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10369_ sha256cu.msg_scheduler.mreg_6\[1\] _04434_ _04446_ _04437_ VGND VGND VPWR
+ VPWR _00653_ sky130_fd_sc_hd__o211a_1
X_13157_ _06573_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__clkbuf_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ sha256cu.msg_scheduler.mreg_1\[25\] sha256cu.msg_scheduler.mreg_1\[8\] VGND
+ VGND VPWR VPWR _05919_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _06536_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__clkbuf_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12039_ _05850_ _05851_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__and2_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_07580_ _02202_ _02204_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09250_ _03729_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__nand2_1
X_08201_ sha256cu.m_out_digest.h_in\[22\] _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__xnor2_1
X_09181_ _03606_ _03636_ _03635_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__a21oi_1
XFILLER_146_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08132_ sha256cu.iter_processing.w\[20\] _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__xor2_2
XFILLER_134_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08063_ sha256cu.m_out_digest.e_in\[29\] _02674_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__xnor2_4
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07014_ _01617_ _01614_ _01695_ _01697_ _01698_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__a32o_1
XFILLER_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08965_ _02380_ _03423_ _03424_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__a21boi_1
XFILLER_115_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput208 hash[56] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
X_07916_ _02493_ _02496_ _02531_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__o21a_1
XFILLER_57_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput219 hash[66] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_4
X_08896_ _03336_ _03361_ _03360_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__a21o_1
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07847_ _02410_ _02429_ _02464_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__a21bo_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07778_ sha256cu.K\[10\] _02397_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09517_ _03082_ _03959_ _03958_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__a21boi_1
XFILLER_72_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _03890_ _03894_ _03921_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__a21oi_1
XFILLER_40_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09379_ _03850_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nor2_1
XFILLER_8_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12390_ _06164_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__clkbuf_1
X_11410_ _05125_ _05139_ _05232_ _05241_ _05253_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__a311o_1
XFILLER_137_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11341_ _05182_ _05184_ _05189_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__or3_1
XFILLER_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14060_ clknet_leaf_39_clk _00606_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11272_ sha256cu.data_in_padd\[15\] _01963_ _05094_ _05123_ _05040_ VGND VGND VPWR
+ VPWR _00878_ sky130_fd_sc_hd__o221a_1
XFILLER_4_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10223_ sha256cu.msg_scheduler.mreg_4\[2\] _04354_ _04363_ _04357_ VGND VGND VPWR
+ VPWR _00590_ sky130_fd_sc_hd__o211a_1
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13011_ _06495_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10154_ sha256cu.msg_scheduler.mreg_3\[4\] _04315_ _04324_ _04318_ VGND VGND VPWR
+ VPWR _00560_ sky130_fd_sc_hd__o211a_1
XFILLER_121_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10085_ sha256cu.msg_scheduler.mreg_3\[7\] _04282_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__or2_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14893_ clknet_leaf_10_clk _01407_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13913_ clknet_leaf_105_clk _00459_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.temp_case
+ sky130_fd_sc_hd__dfxtp_1
X_13844_ clknet_leaf_17_clk _00390_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13775_ clknet_leaf_73_clk _00321_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10987_ sha256cu.m_pad_pars.block_512\[15\]\[2\] _04781_ _04851_ _01970_ VGND VGND
+ VPWR VPWR _04852_ sky130_fd_sc_hd__a211o_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12726_ sha256cu.m_pad_pars.block_512\[22\]\[0\] _06343_ VGND VGND VPWR VPWR _06344_
+ sky130_fd_sc_hd__and2_1
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12657_ _06251_ _05081_ _04994_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__or3_4
XFILLER_31_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11608_ sha256cu.msg_scheduler.mreg_14\[19\] _05440_ VGND VGND VPWR VPWR _05441_
+ sky130_fd_sc_hd__xnor2_1
X_12588_ _01964_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__buf_6
X_14327_ clknet_leaf_89_clk _00021_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11539_ sha256cu.m_pad_pars.block_512\[8\]\[6\] _05318_ _05299_ sha256cu.m_pad_pars.block_512\[12\]\[6\]
+ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__a22o_1
XFILLER_144_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14258_ clknet_leaf_25_clk _00804_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_14189_ clknet_leaf_29_clk _00735_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13209_ _06601_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _02081_ _03227_ _03226_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__a21boi_1
XFILLER_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07701_ _02320_ _02322_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__xor2_2
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08681_ sha256cu.m_out_digest.d_in\[23\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[23\]
+ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__a22o_1
X_07632_ _02252_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__or2_1
XFILLER_93_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07563_ sha256cu.m_out_digest.b_in\[5\] sha256cu.m_out_digest.a_in\[5\] VGND VGND
+ VPWR VPWR _02188_ sky130_fd_sc_hd__or2_1
X_09302_ _03717_ _03750_ _03749_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a21oi_2
XFILLER_53_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07494_ _02118_ _02119_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__and3_1
XFILLER_22_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09233_ _03713_ _03714_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__xor2_1
X_09164_ _02643_ _03617_ _03618_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__a21boi_1
X_08115_ _02703_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__xor2_2
XFILLER_119_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09095_ _03551_ _03557_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__and3_1
XFILLER_108_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08046_ _02632_ _02617_ _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__and3_1
XFILLER_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09997_ _04166_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__buf_2
XFILLER_130_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08948_ _03438_ _03439_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__xnor2_1
X_08879_ _02270_ _03349_ _03350_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__a21bo_1
XFILLER_57_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10910_ _04748_ _04776_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__nor2_2
X_11890_ sha256cu.iter_processing.w\[12\] _05666_ _05710_ _05640_ VGND VGND VPWR VPWR
+ _00910_ sky130_fd_sc_hd__o211a_1
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10841_ sha256cu.m_pad_pars.add_out2\[2\] _01963_ _01966_ VGND VGND VPWR VPWR _04719_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10772_ sha256cu.msg_scheduler.mreg_11\[14\] _04672_ _04676_ _04675_ VGND VGND VPWR
+ VPWR _00826_ sky130_fd_sc_hd__o211a_1
X_13560_ clknet_leaf_68_clk _00106_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[11\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13491_ _06730_ _06758_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__and2_1
X_12511_ _06228_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12442_ sha256cu.m_pad_pars.block_512\[5\]\[4\] _06187_ VGND VGND VPWR VPWR _06192_
+ sky130_fd_sc_hd__and2_1
XFILLER_138_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12373_ sha256cu.m_pad_pars.block_512\[1\]\[3\] _06152_ VGND VGND VPWR VPWR _06156_
+ sky130_fd_sc_hd__and2_1
X_14112_ clknet_leaf_36_clk _00658_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11324_ sha256cu.m_pad_pars.block_512\[29\]\[1\] _05141_ _05138_ sha256cu.m_pad_pars.block_512\[17\]\[1\]
+ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__a221o_1
XFILLER_153_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14043_ clknet_leaf_42_clk _00589_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11255_ _04759_ _04807_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__nor2_1
XFILLER_140_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10206_ sha256cu.msg_scheduler.mreg_3\[27\] _04341_ _04353_ _04344_ VGND VGND VPWR
+ VPWR _00583_ sky130_fd_sc_hd__o211a_1
XFILLER_122_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11186_ sha256cu.m_pad_pars.block_512\[62\]\[3\] _04984_ _04982_ sha256cu.m_pad_pars.block_512\[58\]\[3\]
+ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__a22o_1
X_10137_ _04043_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__buf_2
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10068_ sha256cu.msg_scheduler.mreg_3\[0\] _04268_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__or2_1
X_14945_ clknet_leaf_91_clk _01459_ VGND VGND VPWR VPWR sha256cu.K\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14876_ clknet_leaf_125_clk _01390_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13827_ clknet_leaf_110_clk _00373_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[22\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_63_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13758_ clknet_leaf_70_clk _00304_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12709_ sha256cu.m_pad_pars.block_512\[21\]\[0\] _06334_ VGND VGND VPWR VPWR _06335_
+ sky130_fd_sc_hd__and2_1
X_13689_ clknet_leaf_64_clk _00235_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_117_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09920_ sha256cu.msg_scheduler.mreg_1\[0\] _04174_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__or2_1
XFILLER_125_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09851_ sha256cu.msg_scheduler.mreg_13\[12\] _04147_ VGND VGND VPWR VPWR _04149_
+ sky130_fd_sc_hd__or2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _03297_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__or2b_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09782_ sha256cu.msg_scheduler.mreg_14\[15\] _04106_ VGND VGND VPWR VPWR _04109_
+ sky130_fd_sc_hd__or2_1
XFILLER_39_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06994_ _00454_ _01637_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__nand2_1
XFILLER_105_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08733_ _03208_ _03209_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__or2_1
XFILLER_39_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08664_ sha256cu.m_out_digest.d_in\[8\] _03187_ _03186_ sha256cu.m_out_digest.c_in\[8\]
+ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__o22a_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07615_ _02197_ _02201_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__o21a_1
X_08595_ sha256cu.m_out_digest.b_in\[16\] _02370_ _03176_ _02128_ VGND VGND VPWR VPWR
+ _00143_ sky130_fd_sc_hd__o22a_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _02124_ _02135_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__o21ba_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07477_ _02101_ _02103_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__nor2_1
X_09216_ _03696_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__nand2_1
X_09147_ _03630_ _03631_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__and2_1
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09078_ _02526_ _03535_ _03534_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__o21a_1
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpassword_cracker_264 VGND VGND VPWR VPWR password_cracker_264/HI password_count[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpassword_cracker_286 VGND VGND VPWR VPWR password_cracker_286/HI password_count[26]
+ sky130_fd_sc_hd__conb_1
X_08029_ sha256cu.m_out_digest.e_in\[23\] sha256cu.m_out_digest.e_in\[10\] VGND VGND
+ VPWR VPWR _02642_ sky130_fd_sc_hd__xnor2_2
Xpassword_cracker_275 VGND VGND VPWR VPWR password_cracker_275/HI password_count[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11040_ sha256cu.m_pad_pars.block_512\[7\]\[6\] _04774_ _04822_ sha256cu.m_pad_pars.block_512\[47\]\[6\]
+ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a22o_1
XFILLER_131_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12991_ sha256cu.m_pad_pars.block_512\[37\]\[4\] _06480_ VGND VGND VPWR VPWR _06485_
+ sky130_fd_sc_hd__and2_1
X_11942_ _05757_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__xor2_1
X_14730_ clknet_leaf_7_clk _01244_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[38\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11873_ _05668_ _05672_ _05669_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__a21boi_1
XFILLER_72_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14661_ clknet_leaf_98_clk _01175_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13612_ clknet_leaf_71_clk _00158_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14592_ clknet_leaf_98_clk _01106_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10824_ sha256cu.m_pad_pars.add_512_block\[1\] _04700_ _04708_ _04709_ VGND VGND
+ VPWR VPWR _00845_ sky130_fd_sc_hd__o211a_1
XFILLER_111_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13543_ clknet_leaf_107_clk _00089_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10755_ sha256cu.msg_scheduler.mreg_12\[7\] _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__or2_1
XFILLER_146_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10686_ sha256cu.msg_scheduler.mreg_11\[9\] _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__or2_1
XFILLER_9_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13474_ sha256cu.K\[16\] _06714_ _06719_ _00043_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__a22o_1
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12425_ sha256cu.m_pad_pars.block_512\[4\]\[4\] _06178_ VGND VGND VPWR VPWR _06183_
+ sky130_fd_sc_hd__and2_1
X_12356_ _06147_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ _01985_ _05152_ _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__and3_2
XFILLER_153_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12287_ _06064_ _06068_ _06089_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__nand3_2
XFILLER_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14026_ clknet_leaf_56_clk _00572_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11238_ _04698_ _04785_ _04786_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__and3_1
XFILLER_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11169_ sha256cu.m_pad_pars.block_512\[50\]\[1\] _05008_ _04981_ sha256cu.m_pad_pars.block_512\[54\]\[1\]
+ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__a221o_1
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14928_ clknet_leaf_95_clk _01442_ VGND VGND VPWR VPWR sha256cu.K\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14859_ clknet_leaf_7_clk _01373_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_07400_ sha256cu.m_out_digest.h_in\[0\] _02029_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08380_ sha256cu.K\[26\] _02983_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__and2b_1
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07331_ _01973_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__clkbuf_8
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07262_ sha256cu.m_pad_pars.add_512_block\[2\] sha256cu.m_pad_pars.add_512_block\[1\]
+ sha256cu.m_pad_pars.add_512_block\[0\] sha256cu.m_pad_pars.add_512_block\[3\] VGND
+ VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a31o_1
X_09001_ _03489_ _03490_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__and2_1
X_07193_ _01631_ _01854_ _01855_ _01857_ _01858_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a32o_1
XFILLER_145_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09903_ sha256cu.msg_scheduler.counter_iteration\[2\] _04178_ _04177_ VGND VGND VPWR
+ VPWR _04180_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09834_ sha256cu.msg_scheduler.mreg_13\[5\] _04134_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__or2_1
XFILLER_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09765_ _04044_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__buf_2
XFILLER_55_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06977_ _00452_ _01600_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__or2_2
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08716_ _03202_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__xnor2_1
X_09696_ _04044_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__buf_2
XFILLER_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ sha256cu.m_out_digest.c_in\[27\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[27\]
+ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__o22a_1
XFILLER_54_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08578_ sha256cu.m_out_digest.b_in\[0\] _02370_ _02110_ sha256cu.m_out_digest.a_in\[0\]
+ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__o22a_1
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07529_ _02151_ _02152_ _02153_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__a21o_1
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10540_ sha256cu.msg_scheduler.mreg_8\[10\] _04540_ _04544_ _04543_ VGND VGND VPWR
+ VPWR _00726_ sky130_fd_sc_hd__o211a_1
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10471_ sha256cu.msg_scheduler.mreg_8\[13\] _04494_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__or2_1
XFILLER_108_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _06015_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__or2_1
XFILLER_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13190_ _06591_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12141_ sha256cu.msg_scheduler.mreg_14\[10\] sha256cu.msg_scheduler.mreg_14\[8\]
+ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__xor2_1
X_12072_ _05883_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__and2_1
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11023_ sha256cu.m_pad_pars.block_512\[59\]\[5\] _04829_ _04833_ sha256cu.m_pad_pars.block_512\[55\]\[5\]
+ _04884_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__a221o_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12974_ sha256cu.m_pad_pars.block_512\[36\]\[4\] _06471_ VGND VGND VPWR VPWR _06476_
+ sky130_fd_sc_hd__and2_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11925_ _05740_ _05742_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__or2_1
X_14713_ clknet_leaf_126_clk _01227_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ sha256cu.msg_scheduler.mreg_14\[28\] sha256cu.msg_scheduler.mreg_14\[21\]
+ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__xnor2_1
X_14644_ clknet_leaf_3_clk _01158_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10807_ sha256cu.msg_scheduler.mreg_12\[30\] _04692_ VGND VGND VPWR VPWR _04696_
+ sky130_fd_sc_hd__or2_1
X_11787_ _05610_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__nand2_1
XFILLER_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14575_ clknet_leaf_0_clk _01089_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10738_ sha256cu.msg_scheduler.mreg_12\[0\] _04653_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__or2_1
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13526_ clknet_leaf_124_clk _00076_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13457_ _04188_ _00067_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__and2b_1
X_10669_ sha256cu.msg_scheduler.mreg_11\[2\] _04614_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__or2_1
X_12408_ sha256cu.m_pad_pars.block_512\[3\]\[4\] _06169_ VGND VGND VPWR VPWR _06174_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13388_ _06695_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12339_ sha256cu.m_pad_pars.add_512_block\[2\] _06132_ sha256cu.m_pad_pars.add_512_block\[3\]
+ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__a21o_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14009_ clknet_leaf_42_clk _00555_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_06900_ _01577_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_4
X_07880_ _02493_ _02496_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06831_ net94 net97 net96 net99 VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__or4_2
X_09550_ _04017_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09481_ _03927_ _03928_ _03953_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__and3_1
XFILLER_64_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08501_ _03058_ _03076_ _03100_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__or3b_1
X_08432_ _02879_ _02884_ _02988_ _02989_ _03026_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__a2111o_1
XFILLER_36_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08363_ sha256cu.m_out_digest.h_in\[25\] _02928_ _02966_ VGND VGND VPWR VPWR _02967_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07314_ _01917_ _01957_ sha256cu.iter_processing.padding_done VGND VGND VPWR VPWR
+ _01958_ sky130_fd_sc_hd__o21ai_1
X_08294_ _02896_ _02899_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07245_ _00454_ _01824_ _01783_ _01621_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__a211o_1
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07176_ _01608_ _01581_ _01626_ _01653_ _01580_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__o32a_1
XFILLER_118_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09817_ sha256cu.msg_scheduler.mreg_14\[30\] _04120_ VGND VGND VPWR VPWR _04129_
+ sky130_fd_sc_hd__or2_1
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09748_ _01973_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__buf_2
XFILLER_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _05535_ _05536_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__nand2_1
X_09679_ sha256cu.msg_scheduler.mreg_14\[2\] _04045_ _04049_ _04050_ VGND VGND VPWR
+ VPWR _00353_ sky130_fd_sc_hd__o211a_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _06324_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__clkbuf_1
X_11641_ sha256cu.msg_scheduler.mreg_1\[20\] _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__xnor2_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14360_ clknet_leaf_14_clk _00874_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11572_ _01936_ _01992_ _05407_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__and3_1
X_10523_ sha256cu.msg_scheduler.mreg_9\[3\] _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__or2_1
Xinput19 hash[116] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13311_ sha256cu.m_pad_pars.block_512\[56\]\[2\] _01924_ VGND VGND VPWR VPWR _06655_
+ sky130_fd_sc_hd__and2_1
X_14291_ clknet_leaf_25_clk _00837_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10454_ sha256cu.msg_scheduler.mreg_7\[5\] _04487_ _04495_ _04490_ VGND VGND VPWR
+ VPWR _00689_ sky130_fd_sc_hd__o211a_1
X_13242_ sha256cu.m_pad_pars.block_512\[52\]\[1\] _06617_ VGND VGND VPWR VPWR _06619_
+ sky130_fd_sc_hd__and2_1
X_10385_ sha256cu.msg_scheduler.mreg_6\[7\] _04448_ _04456_ _04451_ VGND VGND VPWR
+ VPWR _00659_ sky130_fd_sc_hd__o211a_1
XFILLER_124_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13173_ sha256cu.m_pad_pars.block_512\[48\]\[1\] _06580_ VGND VGND VPWR VPWR _06582_
+ sky130_fd_sc_hd__and2_1
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12124_ _05885_ _05910_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__and2_1
XFILLER_2_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12055_ sha256cu.msg_scheduler.mreg_9\[20\] sha256cu.msg_scheduler.mreg_0\[20\] VGND
+ VGND VPWR VPWR _05868_ sky130_fd_sc_hd__nand2_1
XFILLER_78_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11006_ _04865_ _04867_ _04868_ _04869_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__or4_2
XFILLER_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12957_ sha256cu.m_pad_pars.block_512\[35\]\[4\] _06462_ VGND VGND VPWR VPWR _06467_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ _05704_ _05707_ _05726_ _05432_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__a31o_1
XANTENNA_260 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12888_ sha256cu.m_pad_pars.block_512\[31\]\[4\] _06425_ VGND VGND VPWR VPWR _06430_
+ sky130_fd_sc_hd__and2_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11839_ _05616_ _05641_ _05660_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__a211o_1
XANTENNA_293 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14627_ clknet_leaf_98_clk _01141_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_282 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_271 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14558_ clknet_leaf_117_clk _01072_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14489_ clknet_leaf_121_clk _01003_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13509_ sha256cu.K\[29\] _06713_ _06718_ _00057_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__a22o_1
X_07030_ _01606_ _01602_ _01706_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__and3_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08981_ _03441_ _03448_ _03471_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07932_ _02481_ _02512_ _02510_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__o21a_1
XFILLER_114_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07863_ _02382_ _02070_ _02477_ _02480_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__a22o_1
XFILLER_69_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09602_ sha256cu.m_out_digest.g_in\[6\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[6\]
+ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__a22o_1
XFILLER_113_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06814_ net152 net155 net154 net158 VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__or4_4
XFILLER_84_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07794_ sha256cu.m_out_digest.g_in\[11\] sha256cu.m_out_digest.f_in\[11\] sha256cu.m_out_digest.e_in\[11\]
+ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__mux2_2
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09533_ _04002_ _04003_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__or2_1
XFILLER_37_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09464_ sha256cu.iter_processing.w\[28\] _03052_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__and2_1
XFILLER_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09395_ sha256cu.m_out_digest.h_in\[26\] sha256cu.m_out_digest.d_in\[26\] VGND VGND
+ VPWR VPWR _03871_ sky130_fd_sc_hd__nand2_1
X_08415_ sha256cu.iter_processing.w\[26\] _02972_ _03017_ VGND VGND VPWR VPWR _03018_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_40_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08346_ _02924_ _02950_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__and2_1
XFILLER_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08277_ _02837_ _02881_ _02882_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07228_ _01631_ _01885_ _01886_ _01888_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__a31o_1
XFILLER_146_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07159_ _00457_ _01826_ _01827_ _01829_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10170_ sha256cu.msg_scheduler.mreg_3\[11\] _04328_ _04333_ _04331_ VGND VGND VPWR
+ VPWR _00567_ sky130_fd_sc_hd__o211a_1
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13860_ clknet_leaf_23_clk _00406_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13791_ clknet_leaf_69_clk _00337_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12811_ _06251_ _05081_ _04754_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__or3_4
X_12742_ _06352_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__clkbuf_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _06315_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11624_ _05454_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__xor2_2
XFILLER_70_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14412_ clknet_leaf_110_clk _00926_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[28\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14343_ clknet_leaf_112_clk _00857_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out3\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_11_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11555_ _05277_ _05388_ _05390_ _05297_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__a22o_1
X_10506_ sha256cu.msg_scheduler.mreg_7\[28\] _04513_ _04524_ _04516_ VGND VGND VPWR
+ VPWR _00712_ sky130_fd_sc_hd__o211a_1
X_14274_ clknet_leaf_20_clk _00820_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11486_ sha256cu.m_pad_pars.block_512\[24\]\[1\] _05279_ _05294_ sha256cu.m_pad_pars.block_512\[20\]\[1\]
+ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__a22o_1
X_10437_ sha256cu.msg_scheduler.mreg_6\[30\] _04474_ _04485_ _04477_ VGND VGND VPWR
+ VPWR _00682_ sky130_fd_sc_hd__o211a_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13225_ sha256cu.m_pad_pars.block_512\[51\]\[1\] _06608_ VGND VGND VPWR VPWR _06610_
+ sky130_fd_sc_hd__and2_1
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10368_ sha256cu.msg_scheduler.mreg_7\[1\] _04441_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__or2_1
XFILLER_124_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13156_ sha256cu.m_pad_pars.block_512\[47\]\[1\] _06571_ VGND VGND VPWR VPWR _06573_
+ sky130_fd_sc_hd__and2_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10299_ sha256cu.msg_scheduler.mreg_5\[3\] _04393_ _04406_ _04397_ VGND VGND VPWR
+ VPWR _00623_ sky130_fd_sc_hd__o211a_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12107_ _05916_ _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__nand2_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ sha256cu.m_pad_pars.block_512\[43\]\[1\] _06534_ VGND VGND VPWR VPWR _06536_
+ sky130_fd_sc_hd__and2_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12038_ _05850_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__nor2_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13989_ clknet_leaf_58_clk _00535_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08200_ _02083_ _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__xnor2_1
X_09180_ _03662_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__nor2_1
X_08131_ _02739_ _02740_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__xnor2_2
XFILLER_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08062_ sha256cu.m_out_digest.e_in\[24\] sha256cu.m_out_digest.e_in\[11\] VGND VGND
+ VPWR VPWR _02674_ sky130_fd_sc_hd__xnor2_2
XFILLER_146_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07013_ _01691_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__inv_2
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08964_ _02417_ _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__xnor2_1
Xinput209 hash[57] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07915_ sha256cu.m_out_digest.h_in\[13\] _02495_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__nand2_1
XFILLER_69_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08895_ _03387_ _03388_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__nor2_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07846_ _02428_ _02426_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__or2b_1
XFILLER_110_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07777_ _02394_ _02396_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09516_ _03119_ _03987_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _03890_ _03894_ _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__and3_1
XFILLER_25_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09378_ sha256cu.K\[25\] _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08329_ sha256cu.m_out_digest.h_in\[24\] _02892_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__and2_1
XFILLER_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11340_ sha256cu.m_pad_pars.block_512\[9\]\[2\] _05144_ _05147_ sha256cu.m_pad_pars.block_512\[33\]\[2\]
+ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a221o_1
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13010_ sha256cu.m_pad_pars.block_512\[38\]\[5\] _06489_ VGND VGND VPWR VPWR _06495_
+ sky130_fd_sc_hd__and2_1
X_11271_ _05098_ _05100_ _05116_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__or4b_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10222_ sha256cu.msg_scheduler.mreg_5\[2\] _04361_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__or2_1
XFILLER_4_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10153_ sha256cu.msg_scheduler.mreg_4\[4\] _04322_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__or2_1
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10084_ sha256cu.msg_scheduler.mreg_2\[6\] _04274_ _04284_ _04277_ VGND VGND VPWR
+ VPWR _00530_ sky130_fd_sc_hd__o211a_1
XFILLER_48_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14892_ clknet_leaf_9_clk _01406_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13912_ clknet_leaf_105_clk _00458_ VGND VGND VPWR VPWR sha256cu.counter_iteration\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_13843_ clknet_leaf_17_clk _00389_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13774_ clknet_leaf_71_clk _00320_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10986_ sha256cu.m_pad_pars.block_512\[3\]\[2\] _04765_ _04774_ sha256cu.m_pad_pars.block_512\[7\]\[2\]
+ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a22o_1
XFILLER_16_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12725_ _05011_ _05012_ _06270_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__o21ai_4
XFILLER_15_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12656_ _06306_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__clkbuf_1
X_11607_ sha256cu.msg_scheduler.mreg_14\[17\] sha256cu.msg_scheduler.mreg_14\[10\]
+ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__xnor2_1
X_12587_ _06269_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14326_ clknet_leaf_95_clk _00020_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11538_ sha256cu.data_in_padd\[29\] _01980_ _01987_ _05375_ VGND VGND VPWR VPWR _00892_
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14257_ clknet_leaf_25_clk _00803_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11469_ _04701_ _04768_ _05154_ _01943_ _04761_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__o32a_1
X_14188_ clknet_leaf_29_clk _00734_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_13208_ sha256cu.m_pad_pars.block_512\[50\]\[1\] _06599_ VGND VGND VPWR VPWR _06601_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13139_ sha256cu.m_pad_pars.block_512\[46\]\[1\] _06562_ VGND VGND VPWR VPWR _06564_
+ sky130_fd_sc_hd__and2_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ sha256cu.K\[7\] _02288_ _02321_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__a21o_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08680_ sha256cu.m_out_digest.d_in\[22\] _03191_ _03190_ sha256cu.m_out_digest.c_in\[22\]
+ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__o22a_1
X_07631_ _02183_ _02253_ _02254_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__a21o_1
XFILLER_26_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07562_ sha256cu.iter_processing.w\[4\] _02155_ _02154_ VGND VGND VPWR VPWR _02187_
+ sky130_fd_sc_hd__a21o_1
XFILLER_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09301_ _03725_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07493_ sha256cu.m_out_digest.g_in\[3\] sha256cu.m_out_digest.f_in\[3\] sha256cu.m_out_digest.e_in\[3\]
+ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_62_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09232_ sha256cu.K\[19\] _03677_ _03678_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__a21bo_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09163_ _02675_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__xor2_1
XFILLER_119_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08114_ _02705_ _02724_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09094_ _03579_ _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__nor2_1
X_08045_ sha256cu.K\[17\] _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09996_ sha256cu.msg_scheduler.mreg_1\[1\] _04221_ _04233_ _04224_ VGND VGND VPWR
+ VPWR _00493_ sky130_fd_sc_hd__o211a_1
XFILLER_103_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08947_ sha256cu.K\[9\] _03404_ _03405_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__a21bo_1
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08878_ _02302_ _03371_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__xor2_1
XFILLER_57_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07829_ _02445_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10840_ sha256cu.m_pad_pars.add_out2\[2\] _01961_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__and2_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10771_ sha256cu.msg_scheduler.mreg_12\[14\] _04666_ VGND VGND VPWR VPWR _04676_
+ sky130_fd_sc_hd__or2_1
XFILLER_40_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13490_ sha256cu.K\[22\] _06713_ _06718_ _00050_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__a22o_1
X_12510_ sha256cu.m_pad_pars.block_512\[9\]\[4\] _06223_ VGND VGND VPWR VPWR _06228_
+ sky130_fd_sc_hd__and2_1
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12441_ _06191_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12372_ _06155_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__clkbuf_1
X_14111_ clknet_leaf_36_clk _00657_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11323_ sha256cu.m_pad_pars.block_512\[1\]\[1\] _05135_ _05151_ sha256cu.m_pad_pars.block_512\[49\]\[1\]
+ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_14042_ clknet_leaf_44_clk _00588_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_4\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11254_ _04978_ _05104_ _05105_ _01921_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__a22o_1
XFILLER_4_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10205_ sha256cu.msg_scheduler.mreg_4\[27\] _04348_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__or2_1
X_11185_ sha256cu.m_pad_pars.block_512\[30\]\[3\] _05009_ _04977_ sha256cu.m_pad_pars.block_512\[46\]\[3\]
+ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__a22o_1
X_10136_ sha256cu.msg_scheduler.mreg_2\[29\] _04301_ _04313_ _04304_ VGND VGND VPWR
+ VPWR _00553_ sky130_fd_sc_hd__o211a_1
XFILLER_122_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10067_ _04166_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14944_ clknet_leaf_91_clk _01458_ VGND VGND VPWR VPWR sha256cu.K\[17\] sky130_fd_sc_hd__dfxtp_2
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14875_ clknet_leaf_125_clk _01389_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13826_ clknet_leaf_110_clk _00372_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[21\]
+ sky130_fd_sc_hd__dfxtp_2
X_13757_ clknet_leaf_68_clk _00303_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10969_ sha256cu.m_pad_pars.block_512\[51\]\[0\] _04826_ _04828_ sha256cu.m_pad_pars.block_512\[23\]\[0\]
+ _04835_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__a221o_1
XFILLER_149_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12708_ _06270_ _05156_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__nand2_2
XFILLER_31_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13688_ clknet_leaf_65_clk _00234_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_129_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12639_ _06297_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_1
X_14309_ clknet_leaf_92_clk _00002_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09850_ sha256cu.msg_scheduler.mreg_12\[11\] _04140_ _04148_ _04144_ VGND VGND VPWR
+ VPWR _00426_ sky130_fd_sc_hd__o211a_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08801_ sha256cu.iter_processing.w\[5\] _02190_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__or2_1
XFILLER_100_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09781_ sha256cu.msg_scheduler.mreg_13\[14\] _04099_ _04108_ _04103_ VGND VGND VPWR
+ VPWR _00397_ sky130_fd_sc_hd__o211a_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _01603_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_4
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _03225_ _03231_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__xor2_1
XFILLER_39_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ sha256cu.m_out_digest.d_in\[7\] _03189_ _03188_ sha256cu.m_out_digest.c_in\[7\]
+ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__a22o_1
XFILLER_66_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07614_ sha256cu.m_out_digest.h_in\[5\] _02200_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__nand2_1
X_08594_ _02109_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__buf_4
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07545_ _02132_ _02134_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nor2_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07476_ _02101_ _02103_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__and2_1
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09215_ sha256cu.m_out_digest.h_in\[20\] sha256cu.m_out_digest.d_in\[20\] VGND VGND
+ VPWR VPWR _03697_ sky130_fd_sc_hd__nand2_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09146_ _03590_ _03597_ _03629_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__or3_1
XFILLER_108_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09077_ _02565_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__xor2_1
XFILLER_151_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpassword_cracker_265 VGND VGND VPWR VPWR password_cracker_265/HI password_count[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpassword_cracker_276 VGND VGND VPWR VPWR password_cracker_276/HI password_count[16]
+ sky130_fd_sc_hd__conb_1
X_08028_ sha256cu.iter_processing.w\[17\] _02640_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__xnor2_1
Xpassword_cracker_287 VGND VGND VPWR VPWR password_cracker_287/HI password_count[27]
+ sky130_fd_sc_hd__conb_1
XFILLER_89_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09979_ sha256cu.msg_scheduler.mreg_0\[25\] _04221_ _04223_ _04224_ VGND VGND VPWR
+ VPWR _00485_ sky130_fd_sc_hd__o211a_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12990_ _06484_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__clkbuf_1
X_11941_ sha256cu.msg_scheduler.mreg_1\[22\] _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11872_ _05690_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__xor2_1
XFILLER_55_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14660_ clknet_leaf_98_clk _01174_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[29\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13611_ clknet_leaf_74_clk _00157_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10823_ _01994_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_118_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_16
X_14591_ clknet_leaf_98_clk _01105_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[21\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13542_ clknet_leaf_117_clk _00088_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out0\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_10754_ _04547_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__clkbuf_2
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10685_ _04547_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__clkbuf_2
X_13473_ _06747_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__clkbuf_1
X_12424_ _06182_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12355_ sha256cu.m_pad_pars.block_512\[0\]\[2\] _06144_ VGND VGND VPWR VPWR _06147_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11306_ _05156_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__inv_1
XFILLER_141_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12286_ _06064_ _06068_ _06089_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__a21oi_2
XFILLER_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14025_ clknet_leaf_56_clk _00571_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11237_ _04951_ _04967_ _05085_ _05088_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__a31o_1
XFILLER_95_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11168_ sha256cu.m_pad_pars.block_512\[58\]\[1\] _01921_ _04982_ _05025_ _04984_
+ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__a32o_1
X_10119_ sha256cu.msg_scheduler.mreg_2\[21\] _04301_ _04303_ _04304_ VGND VGND VPWR
+ VPWR _00545_ sky130_fd_sc_hd__o211a_1
XFILLER_121_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11099_ sha256cu.m_pad_pars.add_out2\[2\] sha256cu.m_pad_pars.add_out2\[3\] VGND
+ VGND VPWR VPWR _04958_ sky130_fd_sc_hd__and2b_1
XFILLER_63_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14927_ clknet_leaf_90_clk _01441_ VGND VGND VPWR VPWR sha256cu.K\[0\] sky130_fd_sc_hd__dfxtp_2
X_14858_ clknet_leaf_7_clk _01372_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13809_ clknet_leaf_47_clk _00355_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_109_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_16
X_14789_ clknet_leaf_106_clk _01303_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_07330_ _01972_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__buf_4
XFILLER_149_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09000_ _03475_ _03462_ _03488_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__or3_1
X_07261_ sha256cu.m_pad_pars.add_512_block\[5\] sha256cu.m_pad_pars.add_512_block\[4\]
+ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__and2_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07192_ _01618_ _01748_ _01744_ _01629_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__a31oi_1
XFILLER_145_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09902_ sha256cu.msg_scheduler.counter_iteration\[1\] _04176_ _04179_ VGND VGND VPWR
+ VPWR _00447_ sky130_fd_sc_hd__o21a_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09833_ sha256cu.msg_scheduler.mreg_12\[4\] _04126_ _04138_ _04130_ VGND VGND VPWR
+ VPWR _00419_ sky130_fd_sc_hd__o211a_1
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09764_ sha256cu.msg_scheduler.mreg_13\[7\] _04086_ _04098_ _04090_ VGND VGND VPWR
+ VPWR _00390_ sky130_fd_sc_hd__o211a_1
XFILLER_74_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06976_ _01631_ _01645_ _01651_ _01664_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__o31ai_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ sha256cu.msg_scheduler.mreg_14\[9\] _04045_ _04059_ _04050_ VGND VGND VPWR
+ VPWR _00360_ sky130_fd_sc_hd__o211a_1
X_08715_ _03210_ _03215_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__xor2_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08646_ sha256cu.m_out_digest.c_in\[26\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[26\]
+ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__o22a_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08577_ _02040_ _03173_ _03174_ _03175_ _01984_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__o311a_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07528_ _02151_ _02152_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__and3_1
X_07459_ sha256cu.m_out_digest.h_in\[2\] _02086_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__xnor2_1
X_10470_ sha256cu.msg_scheduler.mreg_7\[12\] _04500_ _04504_ _04503_ VGND VGND VPWR
+ VPWR _00696_ sky130_fd_sc_hd__o211a_1
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09129_ _02040_ _03613_ _03614_ _03366_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__o211a_1
XFILLER_135_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12140_ _05948_ _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__nor2_1
XFILLER_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12071_ _05881_ _05882_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__nand2_1
XFILLER_104_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11022_ sha256cu.m_pad_pars.block_512\[31\]\[5\] _04811_ _04883_ _04738_ VGND VGND
+ VPWR VPWR _04884_ sky130_fd_sc_hd__a22o_1
XFILLER_104_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12973_ _06475_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__clkbuf_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _05740_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__nand2_1
X_14712_ clknet_leaf_125_clk _01226_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ clknet_leaf_3_clk _01157_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _05675_ _05676_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__nor2_1
X_11786_ _05607_ _05609_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__or2_1
X_10806_ sha256cu.msg_scheduler.mreg_11\[29\] _04685_ _04695_ _04688_ VGND VGND VPWR
+ VPWR _00841_ sky130_fd_sc_hd__o211a_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14574_ clknet_leaf_112_clk _01088_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10737_ sha256cu.msg_scheduler.mreg_10\[31\] _04646_ _04656_ _04649_ VGND VGND VPWR
+ VPWR _00811_ sky130_fd_sc_hd__o211a_1
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13525_ clknet_leaf_2_clk _00075_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13456_ sha256cu.K\[8\] _06726_ _06727_ _06736_ _06737_ VGND VGND VPWR VPWR _01449_
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10668_ sha256cu.msg_scheduler.mreg_10\[1\] _04607_ _04617_ _04610_ VGND VGND VPWR
+ VPWR _00781_ sky130_fd_sc_hd__o211a_1
X_12407_ _06173_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10599_ sha256cu.msg_scheduler.mreg_10\[4\] _04574_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__or2_1
X_13387_ sha256cu.m_pad_pars.block_512\[60\]\[6\] _06693_ VGND VGND VPWR VPWR _06695_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12338_ _01947_ _04777_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__and2_1
X_12269_ _06072_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__or2_1
X_14008_ clknet_leaf_41_clk _00554_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06830_ net98 net102 net101 net104 VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__or4_4
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09480_ _03927_ _03928_ _03953_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__a21o_1
X_08500_ _03058_ _03076_ _03100_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__o21ba_1
XFILLER_52_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08431_ _03027_ _03025_ _03032_ _02992_ _03024_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__a221oi_2
XFILLER_51_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08362_ _02929_ _02931_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__and2b_1
XFILLER_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08293_ _02897_ _02851_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__a21oi_1
X_07313_ _01942_ _01944_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07244_ _00455_ _01680_ _01798_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__a21o_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07175_ _01591_ _01666_ _01787_ _01585_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__a211o_1
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09816_ sha256cu.msg_scheduler.mreg_13\[29\] _04126_ _04128_ _04117_ VGND VGND VPWR
+ VPWR _00412_ sky130_fd_sc_hd__o211a_1
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09747_ sha256cu.msg_scheduler.mreg_14\[0\] _04080_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__or2_1
X_06959_ _01608_ _01648_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__nor2_2
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _01973_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__buf_2
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08629_ sha256cu.m_out_digest.c_in\[12\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[12\]
+ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__o22a_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ sha256cu.msg_scheduler.mreg_1\[9\] sha256cu.msg_scheduler.mreg_1\[5\] VGND
+ VGND VPWR VPWR _05471_ sky130_fd_sc_hd__xnor2_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11571_ _04751_ _04769_ _05406_ sha256cu.m_pad_pars.block_512\[12\]\[7\] VGND VGND
+ VPWR VPWR _05407_ sky130_fd_sc_hd__o22a_1
X_10522_ _04414_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13310_ _06654_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
X_14290_ clknet_leaf_25_clk _00836_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10453_ sha256cu.msg_scheduler.mreg_8\[5\] _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__or2_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13241_ _06618_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__clkbuf_1
X_10384_ sha256cu.msg_scheduler.mreg_7\[7\] _04455_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__or2_1
X_13172_ _06581_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12123_ _05933_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__inv_2
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12054_ sha256cu.msg_scheduler.mreg_9\[20\] sha256cu.msg_scheduler.mreg_0\[20\] VGND
+ VGND VPWR VPWR _05867_ sky130_fd_sc_hd__or2_1
XFILLER_96_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11005_ sha256cu.m_pad_pars.block_512\[15\]\[3\] _04781_ _04800_ sha256cu.m_pad_pars.block_512\[39\]\[3\]
+ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__a22o_1
XFILLER_93_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12956_ _06466_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__clkbuf_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _05704_ _05707_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_261 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_250 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12887_ _06429_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _05634_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__inv_2
XANTENNA_294 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_272 net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_283 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14626_ clknet_leaf_96_clk _01140_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14557_ clknet_leaf_119_clk _01071_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_40_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_119_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11769_ _05506_ _05502_ _05523_ _05545_ _05592_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__a2111o_1
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13508_ _06769_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__clkbuf_1
X_14488_ clknet_leaf_120_clk _01002_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13439_ _06716_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08980_ _03469_ _03470_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__nor2_1
X_07931_ _02546_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__inv_2
X_07862_ _02478_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nor2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09601_ sha256cu.m_out_digest.g_in\[5\] _04032_ _04030_ sha256cu.m_out_digest.f_in\[5\]
+ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__o22a_1
XFILLER_84_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06813_ _01507_ _01508_ _01509_ _01510_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__or4_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07793_ sha256cu.m_out_digest.b_in\[11\] sha256cu.m_out_digest.a_in\[11\] _02411_
+ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__o21ai_2
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09532_ _04002_ _04003_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__nand2_1
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09463_ sha256cu.iter_processing.w\[28\] _03052_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__nor2_1
X_09394_ sha256cu.m_out_digest.h_in\[26\] sha256cu.m_out_digest.d_in\[26\] VGND VGND
+ VPWR VPWR _03870_ sky130_fd_sc_hd__or2_1
XFILLER_52_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08414_ _02970_ _02971_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__and2b_1
XFILLER_24_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08345_ _02948_ _02949_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_31_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08276_ _02871_ _02873_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__and2b_1
X_07227_ _01650_ _01700_ _01711_ _01887_ _01663_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__o311a_1
XFILLER_146_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07158_ _01618_ _01828_ _01629_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__o21a_1
XFILLER_133_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07089_ _01657_ _01611_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nor2_1
XFILLER_87_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12810_ _06388_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__clkbuf_1
X_13790_ clknet_leaf_69_clk _00336_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12741_ sha256cu.m_pad_pars.block_512\[22\]\[7\] _05111_ _06351_ VGND VGND VPWR VPWR
+ _06352_ sky130_fd_sc_hd__mux2_1
XFILLER_55_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12672_ sha256cu.m_pad_pars.block_512\[18\]\[7\] _05108_ _06249_ VGND VGND VPWR VPWR
+ _06315_ sky130_fd_sc_hd__mux2_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _05435_ _05438_ _05434_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__a21boi_1
X_14411_ clknet_leaf_109_clk _00925_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[27\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14342_ clknet_leaf_111_clk _00856_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11554_ _04751_ _04917_ _05389_ sha256cu.m_pad_pars.block_512\[44\]\[7\] VGND VGND
+ VPWR VPWR _05390_ sky130_fd_sc_hd__o22a_1
X_10505_ sha256cu.msg_scheduler.mreg_8\[28\] _04520_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__or2_1
X_14273_ clknet_leaf_20_clk _00819_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11485_ sha256cu.m_pad_pars.block_512\[8\]\[1\] _05318_ _05285_ sha256cu.m_pad_pars.block_512\[16\]\[1\]
+ _05326_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__a221o_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10436_ sha256cu.msg_scheduler.mreg_7\[30\] _04481_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__or2_1
X_13224_ _06609_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10367_ sha256cu.msg_scheduler.mreg_6\[0\] _04434_ _04445_ _04437_ VGND VGND VPWR
+ VPWR _00652_ sky130_fd_sc_hd__o211a_1
XFILLER_112_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13155_ _06572_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__clkbuf_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ sha256cu.msg_scheduler.mreg_6\[3\] _04401_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__or2_1
X_12106_ sha256cu.msg_scheduler.mreg_9\[22\] sha256cu.msg_scheduler.mreg_0\[22\] VGND
+ VGND VPWR VPWR _05917_ sky130_fd_sc_hd__nand2_1
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _06535_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__clkbuf_1
X_12037_ _05821_ _05825_ _05822_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__a21boi_1
XFILLER_78_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_89_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_66_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13988_ clknet_leaf_57_clk _00534_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12939_ _06457_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14609_ clknet_leaf_1_clk _01123_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_08130_ sha256cu.m_out_digest.g_in\[20\] sha256cu.m_out_digest.f_in\[20\] sha256cu.m_out_digest.e_in\[20\]
+ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_13_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_21_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08061_ sha256cu.iter_processing.w\[18\] _02672_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07012_ _01657_ _01639_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__or3_1
XFILLER_143_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08963_ _03452_ _03453_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__nor2_1
XFILLER_102_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07914_ _02526_ _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__xnor2_1
X_08894_ _03356_ _03367_ _03386_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__and3_1
XFILLER_84_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07845_ _02443_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__xnor2_1
X_07776_ _02335_ _02356_ _02395_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__a21bo_1
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09515_ _03985_ _03986_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__nor2_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ _03919_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__nor2_1
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09377_ _03852_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__nor2_1
XFILLER_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08328_ sha256cu.m_out_digest.h_in\[24\] _02892_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__or2_1
X_08259_ _02846_ _02822_ _02865_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__o21ba_1
XFILLER_137_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11270_ _04997_ _05119_ _05121_ _04991_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__o22a_1
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10221_ sha256cu.msg_scheduler.mreg_4\[1\] _04354_ _04362_ _04357_ VGND VGND VPWR
+ VPWR _00589_ sky130_fd_sc_hd__o211a_1
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10152_ sha256cu.msg_scheduler.mreg_3\[3\] _04315_ _04323_ _04318_ VGND VGND VPWR
+ VPWR _00559_ sky130_fd_sc_hd__o211a_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10083_ sha256cu.msg_scheduler.mreg_3\[6\] _04282_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__or2_1
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13911_ clknet_leaf_95_clk _00457_ VGND VGND VPWR VPWR sha256cu.counter_iteration\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14891_ clknet_leaf_9_clk _01405_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13842_ clknet_leaf_18_clk _00388_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13773_ clknet_leaf_70_clk _00319_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10985_ sha256cu.data_in_padd\[1\] _04840_ _04842_ _04850_ _01974_ VGND VGND VPWR
+ VPWR _00864_ sky130_fd_sc_hd__o221a_1
XFILLER_16_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12724_ _06342_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12655_ sha256cu.m_pad_pars.block_512\[17\]\[7\] _05266_ _06249_ VGND VGND VPWR VPWR
+ _06306_ sky130_fd_sc_hd__mux2_1
X_11606_ _05436_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12586_ sha256cu.m_pad_pars.block_512\[13\]\[7\] _05258_ _06249_ VGND VGND VPWR VPWR
+ _06269_ sky130_fd_sc_hd__mux2_1
XFILLER_129_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11537_ _05367_ _05369_ _05374_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__or3_2
X_14325_ clknet_leaf_90_clk _00019_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14256_ clknet_leaf_26_clk _00802_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11468_ sha256cu.m_pad_pars.block_512\[32\]\[0\] _05306_ _05310_ sha256cu.m_pad_pars.block_512\[52\]\[0\]
+ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__a22o_1
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10419_ sha256cu.msg_scheduler.mreg_6\[22\] _04474_ _04475_ _04464_ VGND VGND VPWR
+ VPWR _00674_ sky130_fd_sc_hd__o211a_1
XFILLER_124_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14187_ clknet_leaf_29_clk _00733_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13207_ _06600_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__clkbuf_1
X_11399_ _04907_ _05129_ _05242_ sha256cu.m_pad_pars.block_512\[25\]\[7\] VGND VGND
+ VPWR VPWR _05243_ sky130_fd_sc_hd__o22a_1
XFILLER_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13138_ _06563_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__clkbuf_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13069_ _06526_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_39_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07630_ _02186_ _02214_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__and2_1
X_07561_ sha256cu.K\[4\] _02177_ _02185_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09300_ _03719_ _03751_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__nand2_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07492_ sha256cu.m_out_digest.b_in\[3\] sha256cu.m_out_digest.a_in\[3\] sha256cu.m_out_digest.c_in\[3\]
+ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__a21o_1
XFILLER_62_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09231_ _03711_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__and2_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09162_ _03644_ _03645_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__nand2_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08113_ _02721_ _02723_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09093_ _03546_ _03560_ _03578_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a21oi_1
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08044_ _02634_ _02656_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09995_ sha256cu.msg_scheduler.mreg_2\[1\] _04228_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__or2_1
XFILLER_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08946_ _03436_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08877_ _03369_ _03370_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__nand2_1
XFILLER_57_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07828_ sha256cu.m_out_digest.g_in\[12\] sha256cu.m_out_digest.f_in\[12\] sha256cu.m_out_digest.e_in\[12\]
+ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__mux2_2
XFILLER_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07759_ sha256cu.m_out_digest.e_in\[16\] sha256cu.m_out_digest.e_in\[3\] VGND VGND
+ VPWR VPWR _02379_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10770_ sha256cu.msg_scheduler.mreg_11\[13\] _04672_ _04674_ _04675_ VGND VGND VPWR
+ VPWR _00825_ sky130_fd_sc_hd__o211a_1
XFILLER_53_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09429_ _03902_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__nor2_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12440_ sha256cu.m_pad_pars.block_512\[5\]\[3\] _06187_ VGND VGND VPWR VPWR _06191_
+ sky130_fd_sc_hd__and2_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14110_ clknet_leaf_36_clk _00656_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_6\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12371_ sha256cu.m_pad_pars.block_512\[1\]\[2\] _06152_ VGND VGND VPWR VPWR _06155_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11322_ sha256cu.m_pad_pars.block_512\[13\]\[1\] _05128_ _05132_ sha256cu.m_pad_pars.block_512\[41\]\[1\]
+ _05171_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__a221o_1
XFILLER_153_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14041_ clknet_leaf_44_clk _00587_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11253_ sha256cu.m_pad_pars.block_512\[62\]\[7\] _04984_ _04982_ sha256cu.m_pad_pars.block_512\[58\]\[7\]
+ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__a22o_1
XFILLER_4_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10204_ sha256cu.msg_scheduler.mreg_3\[26\] _04341_ _04352_ _04344_ VGND VGND VPWR
+ VPWR _00582_ sky130_fd_sc_hd__o211a_1
X_11184_ sha256cu.data_in_padd\[10\] _04840_ _05036_ _05039_ _05040_ VGND VGND VPWR
+ VPWR _00873_ sky130_fd_sc_hd__o221a_1
X_10135_ sha256cu.msg_scheduler.mreg_3\[29\] _04308_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__or2_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10066_ sha256cu.msg_scheduler.mreg_1\[31\] _04260_ _04273_ _04264_ VGND VGND VPWR
+ VPWR _00523_ sky130_fd_sc_hd__o211a_1
XFILLER_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14943_ clknet_leaf_91_clk _01457_ VGND VGND VPWR VPWR sha256cu.K\[16\] sky130_fd_sc_hd__dfxtp_2
X_14874_ clknet_leaf_125_clk _01388_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13825_ clknet_leaf_110_clk _00371_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[20\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_63_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13756_ clknet_leaf_68_clk _00302_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10968_ sha256cu.m_pad_pars.block_512\[59\]\[0\] _04829_ _04831_ sha256cu.m_pad_pars.block_512\[19\]\[0\]
+ _04834_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__a221o_1
X_13687_ clknet_leaf_65_clk _00233_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[10\]
+ sky130_fd_sc_hd__dfxtp_4
X_12707_ _06333_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_1
X_10899_ sha256cu.m_pad_pars.add_out3\[5\] sha256cu.m_pad_pars.add_out3\[4\] VGND
+ VGND VPWR VPWR _04766_ sky130_fd_sc_hd__nor2_1
X_12638_ sha256cu.m_pad_pars.block_512\[16\]\[7\] _05413_ _06249_ VGND VGND VPWR VPWR
+ _06297_ sky130_fd_sc_hd__mux2_1
XFILLER_11_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ sha256cu.m_pad_pars.block_512\[12\]\[7\] _05407_ _06249_ VGND VGND VPWR VPWR
+ _06260_ sky130_fd_sc_hd__mux2_1
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14308_ clknet_leaf_90_clk _00001_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__dfxtp_1
X_14239_ clknet_leaf_19_clk _00785_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ sha256cu.iter_processing.w\[5\] _02190_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__and2_1
XFILLER_112_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09780_ sha256cu.msg_scheduler.mreg_14\[14\] _04106_ VGND VGND VPWR VPWR _04108_
+ sky130_fd_sc_hd__or2_1
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _01570_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_4
X_08731_ _03229_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ _02923_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__buf_6
X_07613_ _02231_ _02236_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__xnor2_2
XFILLER_66_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08593_ sha256cu.m_out_digest.b_in\[15\] _02370_ _02110_ _02084_ VGND VGND VPWR VPWR
+ _00142_ sky130_fd_sc_hd__o22a_1
XFILLER_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07544_ _02157_ _02169_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__xor2_1
X_07475_ _02035_ _02063_ _02102_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__o21ai_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09214_ sha256cu.m_out_digest.h_in\[20\] sha256cu.m_out_digest.d_in\[20\] VGND VGND
+ VPWR VPWR _03696_ sky130_fd_sc_hd__or2_1
XFILLER_10_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09145_ _03590_ _03597_ _03629_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__o21ai_1
X_09076_ _03561_ _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__nand2_1
Xpassword_cracker_266 VGND VGND VPWR VPWR password_cracker_266/HI password_count[6]
+ sky130_fd_sc_hd__conb_1
Xpassword_cracker_277 VGND VGND VPWR VPWR password_cracker_277/HI password_count[17]
+ sky130_fd_sc_hd__conb_1
X_08027_ _02638_ _02639_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpassword_cracker_288 VGND VGND VPWR VPWR password_cracker_288/HI password_count[28]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09978_ _04116_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__buf_2
XFILLER_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08929_ _03409_ _03408_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__or2b_1
XFILLER_39_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11940_ sha256cu.msg_scheduler.mreg_1\[18\] sha256cu.msg_scheduler.mreg_1\[1\] VGND
+ VGND VPWR VPWR _05758_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11871_ sha256cu.msg_scheduler.mreg_1\[30\] _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13610_ clknet_leaf_82_clk _00156_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14590_ clknet_leaf_117_clk _01104_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[20\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10822_ sha256cu.m_pad_pars.m_size\[4\] _04706_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__or2_1
X_10753_ sha256cu.msg_scheduler.mreg_11\[6\] _04659_ _04665_ _04662_ VGND VGND VPWR
+ VPWR _00818_ sky130_fd_sc_hd__o211a_1
XFILLER_13_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13541_ clknet_leaf_117_clk _00087_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out0\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10684_ sha256cu.msg_scheduler.mreg_10\[8\] _04620_ _04626_ _04623_ VGND VGND VPWR
+ VPWR _00788_ sky130_fd_sc_hd__o211a_1
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13472_ _06730_ _06746_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__and2_1
X_12423_ sha256cu.m_pad_pars.block_512\[4\]\[3\] _06178_ VGND VGND VPWR VPWR _06182_
+ sky130_fd_sc_hd__and2_1
X_12354_ _06146_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11305_ _04746_ _05154_ _05155_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__o21bai_1
XFILLER_153_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14024_ clknet_leaf_57_clk _00570_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12285_ _06087_ _06088_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__xnor2_2
XFILLER_134_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11236_ _04958_ _04967_ _05087_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__and3_1
XFILLER_122_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11167_ sha256cu.m_pad_pars.m_size\[9\] sha256cu.m_pad_pars.block_512\[62\]\[1\]
+ _05024_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__mux2_1
X_10118_ _04263_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__buf_2
XFILLER_110_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11098_ _04952_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__nor2_4
X_10049_ sha256cu.msg_scheduler.mreg_1\[23\] _04260_ _04262_ _04264_ VGND VGND VPWR
+ VPWR _00515_ sky130_fd_sc_hd__o211a_1
X_14926_ clknet_leaf_10_clk _01440_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14857_ clknet_leaf_7_clk _01371_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13808_ clknet_leaf_49_clk _00354_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_90_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14788_ clknet_leaf_106_clk _01302_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13739_ clknet_leaf_70_clk _00285_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07260_ state\[1\] sha256cu.hashing_done _01910_ net257 _01913_ VGND VGND VPWR VPWR
+ _00071_ sky130_fd_sc_hd__a311oi_1
XFILLER_129_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07191_ _01665_ _01647_ _01626_ _01856_ _01650_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__a311o_1
XFILLER_129_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09901_ _04177_ _04178_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nor2_1
XFILLER_99_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09832_ sha256cu.msg_scheduler.mreg_13\[4\] _04134_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__or2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09763_ sha256cu.msg_scheduler.mreg_14\[7\] _04093_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__or2_1
XFILLER_58_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _03211_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06975_ _00456_ _01656_ _01662_ _01663_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__a211o_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ sha256cu.iter_processing.w\[9\] _04054_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__or2_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08645_ sha256cu.m_out_digest.c_in\[25\] _03184_ _03182_ sha256cu.m_out_digest.b_in\[25\]
+ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__a22o_1
XFILLER_26_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ sha256cu.m_out_digest.a_in\[31\] _02439_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__or2_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07527_ sha256cu.m_out_digest.g_in\[4\] sha256cu.m_out_digest.f_in\[4\] sha256cu.m_out_digest.e_in\[4\]
+ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__mux2_1
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07458_ _02083_ _02085_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07389_ sha256cu.m_out_digest.b_in\[0\] sha256cu.m_out_digest.a_in\[0\] _02018_ VGND
+ VGND VPWR VPWR _02019_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09128_ sha256cu.m_out_digest.e_in\[16\] _02439_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__or2_1
XFILLER_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09059_ _03532_ _03517_ _03545_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__or3_1
XFILLER_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12070_ _05881_ _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__or2_1
XFILLER_89_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11021_ sha256cu.m_pad_pars.m_size\[5\] sha256cu.m_pad_pars.block_512\[63\]\[5\]
+ _01919_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__mux2_1
XFILLER_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12972_ sha256cu.m_pad_pars.block_512\[36\]\[3\] _06471_ VGND VGND VPWR VPWR _06475_
+ sky130_fd_sc_hd__and2_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_410 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11923_ sha256cu.msg_scheduler.mreg_14\[31\] _05741_ VGND VGND VPWR VPWR _05742_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14711_ clknet_leaf_120_clk _01225_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[36\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _05673_ _05674_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__and2_1
X_14642_ clknet_leaf_10_clk _01156_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ sha256cu.msg_scheduler.mreg_12\[29\] _04692_ VGND VGND VPWR VPWR _04695_
+ sky130_fd_sc_hd__or2_1
XFILLER_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11785_ _05607_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nand2_1
X_14573_ clknet_leaf_16_clk _01087_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10736_ sha256cu.msg_scheduler.mreg_11\[31\] _04653_ VGND VGND VPWR VPWR _04656_
+ sky130_fd_sc_hd__or2_1
X_13524_ clknet_leaf_1_clk _00074_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10667_ sha256cu.msg_scheduler.mreg_11\[1\] _04614_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__or2_1
X_13455_ _01973_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__buf_2
XFILLER_127_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12406_ sha256cu.m_pad_pars.block_512\[3\]\[3\] _06169_ VGND VGND VPWR VPWR _06173_
+ sky130_fd_sc_hd__and2_1
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10598_ sha256cu.msg_scheduler.mreg_9\[3\] _04567_ _04577_ _04570_ VGND VGND VPWR
+ VPWR _00751_ sky130_fd_sc_hd__o211a_1
X_13386_ _06694_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12337_ sha256cu.m_pad_pars.add_512_block\[2\] _06132_ _06135_ VGND VGND VPWR VPWR
+ _00932_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12268_ _06070_ _06071_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__and2_1
X_14007_ clknet_leaf_41_clk _00553_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11219_ sha256cu.m_pad_pars.block_512\[6\]\[6\] _04957_ _04989_ sha256cu.m_pad_pars.block_512\[14\]\[6\]
+ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__a221o_1
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12199_ _06005_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__nand2_1
XFILLER_110_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput190 hash[3] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_64_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14909_ clknet_leaf_124_clk _01423_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_08430_ _02988_ _03026_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__nor2_1
XFILLER_17_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08361_ _02962_ _02964_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ sha256cu.m_out_digest.h_in\[23\] _02848_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__and2_1
X_07312_ sha256cu.m_pad_pars.temp_chk VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__clkinv_2
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07243_ _01631_ _01898_ _01899_ _01901_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__a31o_1
XFILLER_118_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07174_ _01631_ _01838_ _01842_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09815_ sha256cu.msg_scheduler.mreg_14\[29\] _04120_ VGND VGND VPWR VPWR _04128_
+ sky130_fd_sc_hd__or2_1
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09746_ sha256cu.msg_scheduler.mreg_14\[31\] _04086_ _04088_ _04077_ VGND VGND VPWR
+ VPWR _00382_ sky130_fd_sc_hd__o211a_1
XFILLER_74_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06958_ _01573_ _01606_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__nand2_4
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ sha256cu.iter_processing.w\[2\] _04046_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__or2_1
XFILLER_55_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08628_ sha256cu.m_out_digest.c_in\[11\] _03179_ _03182_ sha256cu.m_out_digest.b_in\[11\]
+ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__a22o_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _01564_ _01582_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__nand2_4
XFILLER_27_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ sha256cu.m_out_digest.g_in\[31\] sha256cu.m_out_digest.f_in\[31\] sha256cu.m_out_digest.e_in\[31\]
+ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__mux2_1
XFILLER_70_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11570_ _05248_ _04698_ _04786_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__and3b_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10521_ sha256cu.msg_scheduler.mreg_8\[2\] _04526_ _04533_ _04530_ VGND VGND VPWR
+ VPWR _00718_ sky130_fd_sc_hd__o211a_1
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13240_ sha256cu.m_pad_pars.block_512\[52\]\[0\] _06617_ VGND VGND VPWR VPWR _06618_
+ sky130_fd_sc_hd__and2_1
X_10452_ _04414_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__clkbuf_2
XFILLER_108_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10383_ _04414_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__clkbuf_2
XFILLER_136_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13171_ sha256cu.m_pad_pars.block_512\[48\]\[0\] _06580_ VGND VGND VPWR VPWR _06581_
+ sky130_fd_sc_hd__and2_1
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12122_ _05931_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__or2_1
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12053_ sha256cu.iter_processing.w\[19\] _05666_ _05865_ _05866_ VGND VGND VPWR VPWR
+ _00917_ sky130_fd_sc_hd__o211a_1
XFILLER_2_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11004_ sha256cu.m_pad_pars.block_512\[11\]\[3\] _04790_ _04831_ sha256cu.m_pad_pars.block_512\[19\]\[3\]
+ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__a22o_1
XFILLER_133_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12955_ sha256cu.m_pad_pars.block_512\[35\]\[3\] _06462_ VGND VGND VPWR VPWR _06466_
+ sky130_fd_sc_hd__and2_1
XFILLER_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11906_ _05724_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__or2b_1
XFILLER_93_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_240 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_251 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12886_ sha256cu.m_pad_pars.block_512\[31\]\[3\] _06425_ VGND VGND VPWR VPWR _06429_
+ sky130_fd_sc_hd__and2_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _05658_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__nand2_1
XANTENNA_273 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_295 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_262 net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_284 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14625_ clknet_leaf_98_clk _01139_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11768_ _05565_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__or2_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ clknet_leaf_120_clk _01070_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10719_ _04580_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13507_ _01975_ _06768_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__and2_1
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11699_ sha256cu.iter_processing.w\[4\] _04043_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__or2_1
X_14487_ clknet_leaf_120_clk _01001_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13438_ _06725_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__clkbuf_1
X_13369_ _06685_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07930_ _02512_ _02470_ _02510_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__nor3b_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07861_ _02470_ _02476_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__nor2_1
XFILLER_110_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07792_ sha256cu.m_out_digest.b_in\[11\] sha256cu.m_out_digest.a_in\[11\] sha256cu.m_out_digest.c_in\[11\]
+ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a21o_1
X_09600_ sha256cu.m_out_digest.g_in\[4\] _04033_ _04031_ sha256cu.m_out_digest.f_in\[4\]
+ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__a22o_1
XFILLER_110_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06812_ net143 net147 net146 net149 VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__or4_4
X_09531_ _03975_ _03976_ _03973_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__a21o_1
X_09462_ _03934_ _03935_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__or2_1
X_09393_ _03832_ _03864_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__and2_1
XFILLER_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08413_ _03013_ _03015_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__xor2_1
XFILLER_12_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08344_ _02909_ _02911_ _02907_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__o21ba_1
XFILLER_51_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08275_ _02873_ _02871_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__or2b_1
X_07226_ _01620_ _01628_ _01872_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__or3_1
XFILLER_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07157_ _01607_ _01690_ _01766_ _01700_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__a31o_1
XFILLER_3_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07088_ _01766_ _01762_ _01617_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__a21o_1
XFILLER_133_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09729_ sha256cu.iter_processing.w\[24\] _04067_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__or2_1
XFILLER_55_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ _01964_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__buf_4
X_12671_ _06314_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11622_ _05451_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__xor2_2
X_14410_ clknet_leaf_109_clk _00924_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[26\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ clknet_leaf_111_clk _00855_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11553_ _04794_ _05248_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__nor2_1
X_10504_ sha256cu.msg_scheduler.mreg_7\[27\] _04513_ _04523_ _04516_ VGND VGND VPWR
+ VPWR _00711_ sky130_fd_sc_hd__o211a_1
XFILLER_109_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14272_ clknet_leaf_20_clk _00818_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11484_ sha256cu.m_pad_pars.block_512\[36\]\[1\] _05304_ _05325_ _01920_ VGND VGND
+ VPWR VPWR _05326_ sky130_fd_sc_hd__a22o_1
XFILLER_137_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10435_ sha256cu.msg_scheduler.mreg_6\[29\] _04474_ _04484_ _04477_ VGND VGND VPWR
+ VPWR _00681_ sky130_fd_sc_hd__o211a_1
X_13223_ sha256cu.m_pad_pars.block_512\[51\]\[0\] _06608_ VGND VGND VPWR VPWR _06609_
+ sky130_fd_sc_hd__and2_1
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13154_ sha256cu.m_pad_pars.block_512\[47\]\[0\] _06571_ VGND VGND VPWR VPWR _06572_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10366_ sha256cu.msg_scheduler.mreg_7\[0\] _04441_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__or2_1
X_12105_ sha256cu.msg_scheduler.mreg_9\[22\] sha256cu.msg_scheduler.mreg_0\[22\] VGND
+ VGND VPWR VPWR _05916_ sky130_fd_sc_hd__or2_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ sha256cu.msg_scheduler.mreg_5\[2\] _04393_ _04405_ _04397_ VGND VGND VPWR
+ VPWR _00622_ sky130_fd_sc_hd__o211a_1
XFILLER_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ sha256cu.m_pad_pars.block_512\[43\]\[0\] _06534_ VGND VGND VPWR VPWR _06535_
+ sky130_fd_sc_hd__and2_1
X_12036_ _05847_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__xor2_1
XFILLER_19_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13987_ clknet_leaf_57_clk _00533_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12938_ sha256cu.m_pad_pars.block_512\[34\]\[3\] _06453_ VGND VGND VPWR VPWR _06457_
+ sky130_fd_sc_hd__and2_1
XFILLER_74_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ sha256cu.m_pad_pars.block_512\[30\]\[3\] _06416_ VGND VGND VPWR VPWR _06420_
+ sky130_fd_sc_hd__and2_1
X_14608_ clknet_leaf_2_clk _01122_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14539_ clknet_leaf_9_clk _01053_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_08060_ _02670_ _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07011_ _01667_ _01634_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__nor2_2
XFILLER_127_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08962_ sha256cu.m_out_digest.h_in\[11\] sha256cu.m_out_digest.d_in\[11\] VGND VGND
+ VPWR VPWR _03453_ sky130_fd_sc_hd__and2_1
XFILLER_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08893_ _03356_ _03367_ _03386_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__a21oi_1
X_07913_ sha256cu.m_out_digest.h_in\[14\] _02528_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07844_ _02459_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07775_ _02355_ _02353_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__or2b_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09514_ sha256cu.m_out_digest.h_in\[30\] sha256cu.m_out_digest.d_in\[30\] VGND VGND
+ VPWR VPWR _03986_ sky130_fd_sc_hd__and2_1
XFILLER_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09445_ _03883_ _03898_ _03918_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__a21oi_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09376_ sha256cu.iter_processing.w\[25\] _02939_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__and2_1
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08327_ _02929_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08258_ _02862_ _02864_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07209_ _01608_ _01602_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__nor2_1
X_10220_ sha256cu.msg_scheduler.mreg_5\[1\] _04361_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__or2_1
X_08189_ _02796_ _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__nand2_1
XFILLER_106_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10151_ sha256cu.msg_scheduler.mreg_4\[3\] _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__or2_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10082_ sha256cu.msg_scheduler.mreg_2\[5\] _04274_ _04283_ _04277_ VGND VGND VPWR
+ VPWR _00529_ sky130_fd_sc_hd__o211a_1
XFILLER_0_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13910_ clknet_leaf_96_clk _00456_ VGND VGND VPWR VPWR sha256cu.counter_iteration\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14890_ clknet_leaf_9_clk _01404_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[58\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13841_ clknet_leaf_18_clk _00387_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13772_ clknet_leaf_70_clk _00318_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10984_ sha256cu.m_pad_pars.block_512\[31\]\[1\] _04811_ _04845_ _04849_ VGND VGND
+ VPWR VPWR _04850_ sky130_fd_sc_hd__a211o_1
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12723_ sha256cu.m_pad_pars.block_512\[21\]\[7\] _05236_ _06249_ VGND VGND VPWR VPWR
+ _06342_ sky130_fd_sc_hd__mux2_1
XFILLER_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12654_ _06305_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__clkbuf_1
X_11605_ sha256cu.msg_scheduler.mreg_1\[18\] _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12585_ _06268_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11536_ sha256cu.m_pad_pars.block_512\[0\]\[5\] _05314_ _05370_ _05373_ VGND VGND
+ VPWR VPWR _05374_ sky130_fd_sc_hd__a211o_1
X_14324_ clknet_leaf_90_clk _00018_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__dfxtp_1
X_14255_ clknet_leaf_26_clk _00801_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13206_ sha256cu.m_pad_pars.block_512\[50\]\[0\] _06599_ VGND VGND VPWR VPWR _06600_
+ sky130_fd_sc_hd__and2_1
X_11467_ sha256cu.m_pad_pars.add_out0\[5\] sha256cu.m_pad_pars.add_out0\[4\] _05293_
+ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__and4_2
XFILLER_143_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10418_ sha256cu.msg_scheduler.mreg_7\[22\] _04468_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__or2_1
XFILLER_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14186_ clknet_leaf_29_clk _00732_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11398_ _04960_ _05010_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__nor2_1
X_10349_ sha256cu.msg_scheduler.mreg_5\[24\] _04434_ _04435_ _04424_ VGND VGND VPWR
+ VPWR _00644_ sky130_fd_sc_hd__o211a_1
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13137_ sha256cu.m_pad_pars.block_512\[46\]\[0\] _06562_ VGND VGND VPWR VPWR _06563_
+ sky130_fd_sc_hd__and2_1
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13068_ sha256cu.m_pad_pars.block_512\[42\]\[0\] _06525_ VGND VGND VPWR VPWR _06526_
+ sky130_fd_sc_hd__and2_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _05830_ _05832_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__or2_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07560_ _02174_ _02176_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07491_ sha256cu.m_out_digest.b_in\[3\] sha256cu.m_out_digest.a_in\[3\] VGND VGND
+ VPWR VPWR _02118_ sky130_fd_sc_hd__or2_1
X_09230_ _03695_ _03681_ _03710_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__or3_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09161_ sha256cu.m_out_digest.h_in\[18\] sha256cu.m_out_digest.d_in\[18\] VGND VGND
+ VPWR VPWR _03645_ sky130_fd_sc_hd__nand2_1
XFILLER_147_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09092_ _03546_ _03560_ _03578_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__and3_1
XFILLER_108_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08112_ _02680_ _02682_ _02722_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__o21a_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08043_ _02636_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09994_ sha256cu.msg_scheduler.mreg_1\[0\] _04221_ _04232_ _04224_ VGND VGND VPWR
+ VPWR _00492_ sky130_fd_sc_hd__o211a_1
XFILLER_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08945_ _03403_ _03407_ _03401_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__o21ba_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08876_ sha256cu.m_out_digest.h_in\[8\] sha256cu.m_out_digest.d_in\[8\] VGND VGND
+ VPWR VPWR _03370_ sky130_fd_sc_hd__nand2_1
XFILLER_84_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07827_ sha256cu.m_out_digest.b_in\[12\] _02382_ _02444_ VGND VGND VPWR VPWR _02445_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_45_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07758_ sha256cu.iter_processing.w\[10\] _02377_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07689_ _02308_ _02310_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__xnor2_2
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09428_ _02964_ _03870_ _03871_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__a21boi_1
XFILLER_40_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09359_ _03808_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__inv_2
XFILLER_138_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12370_ _06154_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11321_ sha256cu.m_pad_pars.block_512\[45\]\[1\] _05126_ VGND VGND VPWR VPWR _05171_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14040_ clknet_leaf_41_clk _00586_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11252_ sha256cu.m_pad_pars.block_512\[54\]\[7\] _05103_ _04979_ VGND VGND VPWR VPWR
+ _05104_ sky130_fd_sc_hd__o21a_1
X_10203_ sha256cu.msg_scheduler.mreg_4\[26\] _04348_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__or2_1
XFILLER_121_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11183_ _01973_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__buf_4
X_10134_ sha256cu.msg_scheduler.mreg_2\[28\] _04301_ _04312_ _04304_ VGND VGND VPWR
+ VPWR _00552_ sky130_fd_sc_hd__o211a_1
XFILLER_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10065_ sha256cu.msg_scheduler.mreg_2\[31\] _04268_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__or2_1
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14942_ clknet_leaf_91_clk _01456_ VGND VGND VPWR VPWR sha256cu.K\[15\] sky130_fd_sc_hd__dfxtp_4
X_14873_ clknet_leaf_125_clk _01387_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13824_ clknet_leaf_76_clk _00370_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13755_ clknet_leaf_67_clk _00301_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10967_ sha256cu.m_pad_pars.block_512\[63\]\[0\] _01919_ _04738_ _04833_ sha256cu.m_pad_pars.block_512\[55\]\[0\]
+ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__a32o_1
XFILLER_149_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13686_ clknet_leaf_65_clk _00232_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[9\]
+ sky130_fd_sc_hd__dfxtp_4
X_10898_ _04763_ sha256cu.m_pad_pars.add_out3\[4\] _04735_ _04764_ VGND VGND VPWR
+ VPWR _04765_ sky130_fd_sc_hd__and4bb_4
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12706_ sha256cu.m_pad_pars.block_512\[20\]\[7\] _05396_ _06249_ VGND VGND VPWR VPWR
+ _06333_ sky130_fd_sc_hd__mux2_1
X_12637_ _06296_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12568_ _06259_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11519_ sha256cu.m_pad_pars.block_512\[44\]\[4\] _05298_ _05320_ sha256cu.m_pad_pars.block_512\[40\]\[4\]
+ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__a22o_1
X_12499_ sha256cu.m_pad_pars.block_512\[8\]\[7\] _05424_ _01983_ VGND VGND VPWR VPWR
+ _06222_ sky130_fd_sc_hd__mux2_1
X_14307_ clknet_leaf_90_clk _00031_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__dfxtp_1
X_14238_ clknet_leaf_19_clk _00784_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14169_ clknet_leaf_35_clk _00715_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _01678_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08730_ _02051_ _03206_ _03205_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__a21boi_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ sha256cu.m_out_digest.d_in\[6\] _03184_ _03188_ sha256cu.m_out_digest.c_in\[6\]
+ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__a22o_1
X_07612_ sha256cu.m_out_digest.h_in\[6\] _02235_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__xnor2_2
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08592_ sha256cu.m_out_digest.b_in\[14\] _03031_ _02114_ sha256cu.m_out_digest.a_in\[14\]
+ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__a22o_1
X_07543_ _02166_ _02168_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07474_ sha256cu.K\[1\] _02062_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__nand2_1
XFILLER_62_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09213_ _03674_ _03675_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nor2_1
XFILLER_50_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09144_ _03627_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__nor2_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09075_ sha256cu.m_out_digest.h_in\[15\] sha256cu.m_out_digest.d_in\[15\] VGND VGND
+ VPWR VPWR _03562_ sky130_fd_sc_hd__nand2_1
XFILLER_146_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08026_ sha256cu.m_out_digest.g_in\[17\] sha256cu.m_out_digest.f_in\[17\] sha256cu.m_out_digest.e_in\[17\]
+ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__mux2_1
Xpassword_cracker_267 VGND VGND VPWR VPWR password_cracker_267/HI password_count[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_116_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xpassword_cracker_289 VGND VGND VPWR VPWR password_cracker_289/HI password_count[29]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xpassword_cracker_278 VGND VGND VPWR VPWR password_cracker_278/HI password_count[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_115_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09977_ sha256cu.msg_scheduler.mreg_1\[25\] _04215_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__or2_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08928_ _03420_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08859_ _03352_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11870_ sha256cu.msg_scheduler.mreg_1\[19\] sha256cu.msg_scheduler.mreg_1\[15\] VGND
+ VGND VPWR VPWR _05691_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10821_ _01939_ _04700_ _04707_ _04688_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__o211a_1
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10752_ sha256cu.msg_scheduler.mreg_12\[6\] _04653_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__or2_1
X_13540_ clknet_leaf_112_clk _00086_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13471_ sha256cu.K\[15\] _06714_ _06719_ _00042_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__a22o_1
X_10683_ sha256cu.msg_scheduler.mreg_11\[8\] _04614_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__or2_1
XFILLER_71_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12422_ _06181_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12353_ sha256cu.m_pad_pars.block_512\[0\]\[1\] _06144_ VGND VGND VPWR VPWR _06146_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12284_ sha256cu.msg_scheduler.mreg_14\[16\] sha256cu.msg_scheduler.mreg_14\[14\]
+ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__xor2_2
XFILLER_5_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11304_ _04807_ _04969_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__nor2_1
XFILLER_153_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14023_ clknet_leaf_57_clk _00569_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11235_ _04913_ _04960_ _05086_ sha256cu.m_pad_pars.block_512\[42\]\[7\] VGND VGND
+ VPWR VPWR _05087_ sky130_fd_sc_hd__o22a_1
XFILLER_107_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11166_ _01919_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__buf_4
X_10117_ sha256cu.msg_scheduler.mreg_3\[21\] _04295_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__or2_1
XFILLER_122_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11097_ _04769_ _04954_ _04955_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10048_ _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__buf_2
X_14925_ clknet_leaf_10_clk _01439_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14856_ clknet_leaf_9_clk _01370_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13807_ clknet_leaf_49_clk _00353_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14787_ clknet_leaf_107_clk _01301_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11999_ _05792_ _05795_ _05813_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__and3_1
X_13738_ clknet_leaf_83_clk _00284_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13669_ clknet_leaf_88_clk _00215_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07190_ _01622_ _01696_ _01747_ _01611_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__o22a_1
XFILLER_117_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09900_ sha256cu.msg_scheduler.counter_iteration\[0\] sha256cu.msg_scheduler.temp_case
+ sha256cu.msg_scheduler.counter_iteration\[1\] VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__and3_1
XFILLER_125_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09831_ sha256cu.msg_scheduler.mreg_12\[3\] _04126_ _04137_ _04130_ VGND VGND VPWR
+ VPWR _00418_ sky130_fd_sc_hd__o211a_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09762_ sha256cu.msg_scheduler.mreg_13\[6\] _04086_ _04097_ _04090_ VGND VGND VPWR
+ VPWR _00389_ sky130_fd_sc_hd__o211a_1
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _01570_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_4
X_08713_ _03212_ _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__nand2_1
XFILLER_86_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ sha256cu.msg_scheduler.mreg_14\[8\] _04045_ _04058_ _04050_ VGND VGND VPWR
+ VPWR _00359_ sky130_fd_sc_hd__o211a_1
XFILLER_94_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08644_ sha256cu.m_out_digest.c_in\[24\] _03184_ _03182_ sha256cu.m_out_digest.b_in\[24\]
+ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__a22o_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _03142_ _03145_ _03172_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__and3_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07526_ sha256cu.m_out_digest.b_in\[4\] sha256cu.m_out_digest.a_in\[4\] sha256cu.m_out_digest.c_in\[4\]
+ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__a21o_1
XFILLER_81_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07457_ _02084_ sha256cu.m_out_digest.a_in\[4\] VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07388_ sha256cu.m_out_digest.b_in\[0\] sha256cu.m_out_digest.a_in\[0\] sha256cu.m_out_digest.c_in\[0\]
+ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__a21o_1
X_09127_ _03608_ _03612_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09058_ _03532_ _03517_ _03545_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__o21ai_1
XFILLER_108_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08009_ _02553_ _02583_ _02622_ _02548_ _02585_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__a221oi_4
XFILLER_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11020_ _01971_ _04881_ _04882_ _04709_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__o211a_1
XFILLER_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12971_ _06474_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_400 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ sha256cu.msg_scheduler.mreg_14\[24\] sha256cu.msg_scheduler.mreg_14\[1\]
+ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14710_ clknet_leaf_114_clk _01224_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[35\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_411 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ _05673_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__nor2_1
XFILLER_61_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14641_ clknet_leaf_2_clk _01155_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ sha256cu.msg_scheduler.mreg_11\[28\] _04685_ _04694_ _04688_ VGND VGND VPWR
+ VPWR _00840_ sky130_fd_sc_hd__o211a_1
XFILLER_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ sha256cu.msg_scheduler.mreg_14\[27\] _05608_ VGND VGND VPWR VPWR _05609_
+ sky130_fd_sc_hd__xnor2_1
X_14572_ clknet_leaf_22_clk _01086_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10735_ sha256cu.msg_scheduler.mreg_10\[30\] _04646_ _04655_ _04649_ VGND VGND VPWR
+ VPWR _00810_ sky130_fd_sc_hd__o211a_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13523_ clknet_leaf_125_clk _00073_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10666_ sha256cu.msg_scheduler.mreg_10\[0\] _04607_ _04616_ _04610_ VGND VGND VPWR
+ VPWR _00780_ sky130_fd_sc_hd__o211a_1
X_13454_ _04188_ _00066_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__and2b_1
X_12405_ _06172_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__clkbuf_1
X_13385_ sha256cu.m_pad_pars.block_512\[60\]\[5\] _06693_ VGND VGND VPWR VPWR _06694_
+ sky130_fd_sc_hd__and2_1
X_10597_ sha256cu.msg_scheduler.mreg_10\[3\] _04574_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__or2_1
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12336_ sha256cu.m_pad_pars.add_512_block\[2\] _06132_ _03288_ VGND VGND VPWR VPWR
+ _06135_ sky130_fd_sc_hd__o21ai_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12267_ _06070_ _06071_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__nor2_2
X_14006_ clknet_leaf_41_clk _00552_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12198_ _05967_ _05984_ _05981_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__o21ai_1
X_11218_ sha256cu.m_pad_pars.block_512\[2\]\[6\] _04999_ _04972_ sha256cu.m_pad_pars.block_512\[38\]\[6\]
+ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__a22o_1
XFILLER_150_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11149_ _04725_ _04721_ _04990_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__and4_4
XFILLER_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput180 hash[30] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
Xinput191 hash[40] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
X_14908_ clknet_leaf_123_clk _01422_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14839_ clknet_leaf_119_clk _01353_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[52\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_08360_ sha256cu.m_out_digest.e_in\[19\] _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__xnor2_4
XFILLER_63_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07311_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__inv_2
X_08291_ sha256cu.m_out_digest.h_in\[23\] _02848_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__or2_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07242_ _01668_ _01795_ _01900_ _01663_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__o211a_1
XFILLER_118_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07173_ _01570_ _01839_ _01841_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__or3_1
XFILLER_127_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09814_ sha256cu.msg_scheduler.mreg_13\[28\] _04126_ _04127_ _04117_ VGND VGND VPWR
+ VPWR _00411_ sky130_fd_sc_hd__o211a_1
XFILLER_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09745_ sha256cu.iter_processing.w\[31\] _04080_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__or2_1
XFILLER_74_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06957_ _01646_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__clkbuf_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09676_ sha256cu.msg_scheduler.mreg_14\[1\] _04045_ _04048_ _03366_ VGND VGND VPWR
+ VPWR _00352_ sky130_fd_sc_hd__o211a_1
XFILLER_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06888_ sha256cu.counter_iteration\[4\] sha256cu.msg_scheduler.counter_iteration\[4\]
+ _01568_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__mux2_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _02113_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__buf_4
XFILLER_27_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08558_ sha256cu.m_out_digest.e_in\[24\] _03156_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xnor2_2
XFILLER_70_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07509_ _02124_ _02135_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__xor2_1
X_08489_ _03088_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10520_ sha256cu.msg_scheduler.mreg_9\[2\] _04520_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__or2_1
X_10451_ sha256cu.msg_scheduler.mreg_7\[4\] _04487_ _04493_ _04490_ VGND VGND VPWR
+ VPWR _00688_ sky130_fd_sc_hd__o211a_1
XFILLER_109_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10382_ sha256cu.msg_scheduler.mreg_6\[6\] _04448_ _04454_ _04451_ VGND VGND VPWR
+ VPWR _00658_ sky130_fd_sc_hd__o211a_1
XFILLER_108_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13170_ _02111_ _04705_ _05286_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__or3_2
X_12121_ _05929_ _05930_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__and2_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12052_ _01994_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11003_ sha256cu.m_pad_pars.block_512\[23\]\[3\] _04828_ _04818_ sha256cu.m_pad_pars.block_512\[35\]\[3\]
+ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__a221o_1
XFILLER_2_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12954_ _06465_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__clkbuf_1
X_11905_ _05695_ _05700_ _05723_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__a21o_1
XFILLER_46_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_241 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_252 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12885_ _06428_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_263 net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _05656_ _05657_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__nand2_1
XANTENNA_274 _01543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_285 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14624_ clknet_leaf_98_clk _01138_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11767_ _05564_ _05585_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__or2_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14555_ clknet_leaf_119_clk _01069_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10718_ sha256cu.msg_scheduler.mreg_10\[23\] _04633_ _04645_ _04636_ VGND VGND VPWR
+ VPWR _00803_ sky130_fd_sc_hd__o211a_1
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13506_ sha256cu.K\[28\] _06713_ _06718_ _00056_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__a22o_1
XFILLER_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11698_ sha256cu.data_in_padd\[4\] _05448_ _05463_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__a21o_1
X_14486_ clknet_leaf_114_clk _01000_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10649_ sha256cu.msg_scheduler.mreg_9\[25\] _04594_ _04606_ _04597_ VGND VGND VPWR
+ VPWR _00773_ sky130_fd_sc_hd__o211a_1
X_13437_ _03288_ _06724_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__and2_1
XFILLER_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13368_ sha256cu.m_pad_pars.block_512\[59\]\[5\] _06682_ VGND VGND VPWR VPWR _06685_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12319_ sha256cu.msg_scheduler.mreg_9\[31\] sha256cu.msg_scheduler.mreg_1\[6\] VGND
+ VGND VPWR VPWR _06121_ sky130_fd_sc_hd__xor2_1
XFILLER_87_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13299_ sha256cu.m_pad_pars.block_512\[55\]\[4\] _06644_ VGND VGND VPWR VPWR _06649_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07860_ _02108_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__buf_4
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07791_ sha256cu.iter_processing.w\[10\] _02376_ _02375_ VGND VGND VPWR VPWR _02410_
+ sky130_fd_sc_hd__a21o_1
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06811_ net139 net142 net141 net144 VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__or4_1
XFILLER_96_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09530_ _04000_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__xor2_1
X_09461_ _03932_ _03933_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__and2_1
XFILLER_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09392_ _02220_ _03866_ _03867_ _03868_ _01984_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__o311a_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08412_ _02968_ _02973_ _03014_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__a21bo_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08343_ _02945_ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__xnor2_1
X_08274_ _02839_ _02874_ _02842_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__or3b_1
XFILLER_138_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07225_ _01643_ _00455_ _01604_ _01701_ _01621_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__a221o_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07156_ _01578_ _01625_ _01703_ _01790_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__a31o_1
XFILLER_133_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07087_ _01637_ _01591_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__nand2_1
XFILLER_99_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07989_ sha256cu.m_out_digest.h_in\[16\] _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__xnor2_1
X_09728_ sha256cu.msg_scheduler.mreg_14\[23\] _04073_ _04078_ _04077_ VGND VGND VPWR
+ VPWR _00374_ sky130_fd_sc_hd__o211a_1
XFILLER_90_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09659_ sha256cu.m_out_digest.h_in\[23\] _04039_ _02478_ sha256cu.m_out_digest.g_in\[23\]
+ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__o22a_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ sha256cu.m_pad_pars.block_512\[18\]\[6\] _06307_ VGND VGND VPWR VPWR _06314_
+ sky130_fd_sc_hd__and2_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ sha256cu.msg_scheduler.mreg_1\[19\] _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__xnor2_2
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ clknet_leaf_111_clk _00854_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.add_out2\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11552_ _04907_ _04751_ _05387_ sha256cu.m_pad_pars.block_512\[28\]\[7\] VGND VGND
+ VPWR VPWR _05388_ sky130_fd_sc_hd__o22a_1
X_10503_ sha256cu.msg_scheduler.mreg_8\[27\] _04520_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__or2_1
X_14271_ clknet_leaf_19_clk _00817_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11483_ sha256cu.m_pad_pars.block_512\[60\]\[1\] _01998_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[1\]
+ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__a22o_1
XFILLER_137_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10434_ sha256cu.msg_scheduler.mreg_7\[29\] _04481_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__or2_1
X_13222_ _04823_ _04825_ _01972_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__o21ai_4
XFILLER_152_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10365_ sha256cu.msg_scheduler.mreg_5\[31\] _04434_ _04444_ _04437_ VGND VGND VPWR
+ VPWR _00651_ sky130_fd_sc_hd__o211a_1
XFILLER_124_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13153_ _02111_ _04705_ _04820_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__or3_4
XFILLER_151_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12104_ sha256cu.iter_processing.w\[21\] _05894_ _05915_ _05866_ VGND VGND VPWR VPWR
+ _00919_ sky130_fd_sc_hd__o211a_1
XFILLER_3_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10296_ sha256cu.msg_scheduler.mreg_6\[2\] _04401_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__or2_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ _01986_ _04803_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__or2_2
X_12035_ sha256cu.msg_scheduler.mreg_1\[26\] _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13986_ clknet_leaf_56_clk _00532_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12937_ _06456_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _06419_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ sha256cu.msg_scheduler.mreg_9\[10\] sha256cu.msg_scheduler.mreg_0\[10\] VGND
+ VGND VPWR VPWR _05642_ sky130_fd_sc_hd__or2_1
XFILLER_21_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14607_ clknet_leaf_0_clk _01121_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[23\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ sha256cu.m_pad_pars.block_512\[26\]\[2\] _06380_ VGND VGND VPWR VPWR _06383_
+ sky130_fd_sc_hd__and2_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14538_ clknet_leaf_8_clk _01052_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14469_ clknet_leaf_98_clk _00983_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07010_ _01640_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__nand2_1
XFILLER_115_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08961_ sha256cu.m_out_digest.h_in\[11\] sha256cu.m_out_digest.d_in\[11\] VGND VGND
+ VPWR VPWR _03452_ sky130_fd_sc_hd__nor2_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08892_ _03368_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07912_ sha256cu.m_out_digest.a_in\[27\] _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07843_ _02415_ _02425_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__o21ba_1
XFILLER_111_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07774_ _02371_ _02393_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09513_ sha256cu.m_out_digest.h_in\[30\] sha256cu.m_out_digest.d_in\[30\] VGND VGND
+ VPWR VPWR _03985_ sky130_fd_sc_hd__nor2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09444_ _03883_ _03898_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__and3_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09375_ _03851_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__inv_2
XFILLER_138_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08326_ sha256cu.m_out_digest.e_in\[31\] _02930_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__xnor2_4
X_08257_ _02816_ _02823_ _02863_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08188_ sha256cu.K\[21\] _02795_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__nand2_1
X_07208_ _01643_ _01610_ _01647_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07139_ _01585_ _00455_ _01681_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__and3_1
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10150_ _04281_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__clkbuf_2
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10081_ sha256cu.msg_scheduler.mreg_3\[5\] _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__or2_1
XFILLER_0_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13840_ clknet_leaf_18_clk _00386_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_13\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13771_ clknet_leaf_71_clk _00317_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10983_ sha256cu.m_pad_pars.block_512\[35\]\[1\] _04818_ _04846_ _04848_ VGND VGND
+ VPWR VPWR _04849_ sky130_fd_sc_hd__a211o_1
X_12722_ _06341_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12653_ sha256cu.m_pad_pars.block_512\[17\]\[6\] _06298_ VGND VGND VPWR VPWR _06305_
+ sky130_fd_sc_hd__and2_1
X_11604_ sha256cu.msg_scheduler.mreg_1\[7\] sha256cu.msg_scheduler.mreg_1\[3\] VGND
+ VGND VPWR VPWR _05437_ sky130_fd_sc_hd__xnor2_1
X_12584_ sha256cu.m_pad_pars.block_512\[13\]\[6\] _06261_ VGND VGND VPWR VPWR _06268_
+ sky130_fd_sc_hd__and2_1
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11535_ sha256cu.m_pad_pars.block_512\[20\]\[5\] _05294_ _05288_ sha256cu.m_pad_pars.block_512\[48\]\[5\]
+ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__a221o_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14323_ clknet_leaf_95_clk _00017_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14254_ clknet_leaf_25_clk _00800_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_13205_ _06270_ _05006_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__nand2_2
X_11466_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__inv_1
X_10417_ _04447_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__buf_2
X_14185_ clknet_leaf_29_clk _00731_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11397_ _05152_ _05149_ _05235_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__a31o_1
XFILLER_151_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10348_ sha256cu.msg_scheduler.mreg_6\[24\] _04428_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__or2_1
XFILLER_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13136_ _02111_ _04917_ _04975_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__or3_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10279_ sha256cu.msg_scheduler.mreg_5\[27\] _04387_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__or2_1
X_13067_ _01986_ _05000_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__or2_2
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ _05830_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__nand2_1
XFILLER_78_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13969_ clknet_leaf_53_clk _00515_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[23\]
+ sky130_fd_sc_hd__dfxtp_2
X_07490_ sha256cu.iter_processing.w\[2\] _02077_ _02076_ VGND VGND VPWR VPWR _02117_
+ sky130_fd_sc_hd__a21o_1
XFILLER_62_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09160_ sha256cu.m_out_digest.h_in\[18\] sha256cu.m_out_digest.d_in\[18\] VGND VGND
+ VPWR VPWR _03644_ sky130_fd_sc_hd__or2_1
X_09091_ _03576_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__xnor2_1
X_08111_ _02673_ _02683_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__or2_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08042_ _02652_ _02654_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09993_ sha256cu.msg_scheduler.mreg_2\[0\] _04228_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__or2_1
XFILLER_116_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08944_ _03430_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__xor2_2
XFILLER_131_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08875_ sha256cu.m_out_digest.h_in\[8\] sha256cu.m_out_digest.d_in\[8\] VGND VGND
+ VPWR VPWR _03369_ sky130_fd_sc_hd__or2_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07826_ sha256cu.m_out_digest.b_in\[12\] _02382_ sha256cu.m_out_digest.c_in\[12\]
+ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__a21o_1
XFILLER_29_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07757_ _02375_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__and2b_1
XFILLER_71_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07688_ _02271_ _02276_ _02309_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__o21a_1
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09427_ _03001_ _03901_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__xor2_1
X_09358_ _03782_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__inv_2
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08309_ _02912_ _02913_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__nand2_1
XFILLER_153_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11320_ sha256cu.data_in_padd\[16\] _04741_ _04742_ _05170_ VGND VGND VPWR VPWR _00879_
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09289_ _03764_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__nor2_1
XFILLER_114_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11251_ _04796_ _04824_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__nor2_1
X_10202_ sha256cu.msg_scheduler.mreg_3\[25\] _04341_ _04351_ _04344_ VGND VGND VPWR
+ VPWR _00581_ sky130_fd_sc_hd__o211a_1
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11182_ sha256cu.m_pad_pars.block_512\[22\]\[2\] _05013_ _05038_ _01971_ VGND VGND
+ VPWR VPWR _05039_ sky130_fd_sc_hd__a211o_1
X_10133_ sha256cu.msg_scheduler.mreg_3\[28\] _04308_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__or2_1
XFILLER_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10064_ sha256cu.msg_scheduler.mreg_1\[30\] _04260_ _04272_ _04264_ VGND VGND VPWR
+ VPWR _00522_ sky130_fd_sc_hd__o211a_1
XFILLER_94_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14941_ clknet_leaf_91_clk _01455_ VGND VGND VPWR VPWR sha256cu.K\[14\] sky130_fd_sc_hd__dfxtp_4
XFILLER_87_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14872_ clknet_leaf_125_clk _01386_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13823_ clknet_leaf_76_clk _00369_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_90_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13754_ clknet_leaf_67_clk _00300_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10966_ _04736_ _04767_ _04832_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__and3_2
X_13685_ clknet_leaf_65_clk _00231_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[8\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_71_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10897_ sha256cu.m_pad_pars.add_out3\[3\] sha256cu.m_pad_pars.add_out3\[2\] VGND
+ VGND VPWR VPWR _04764_ sky130_fd_sc_hd__nor2_2
X_12705_ _06332_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12636_ sha256cu.m_pad_pars.block_512\[16\]\[6\] _06289_ VGND VGND VPWR VPWR _06296_
+ sky130_fd_sc_hd__and2_1
XFILLER_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12567_ sha256cu.m_pad_pars.block_512\[12\]\[6\] _06252_ VGND VGND VPWR VPWR _06259_
+ sky130_fd_sc_hd__and2_1
XFILLER_12_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14306_ clknet_leaf_95_clk _00030_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__dfxtp_1
X_11518_ sha256cu.m_pad_pars.block_512\[32\]\[4\] _05306_ _05318_ sha256cu.m_pad_pars.block_512\[8\]\[4\]
+ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__a221o_1
X_12498_ _06221_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14237_ clknet_leaf_19_clk _00783_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11449_ _04760_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__nor2_1
XFILLER_152_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14168_ clknet_leaf_34_clk _00714_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13119_ _02111_ _04917_ _05124_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__or3_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14099_ clknet_leaf_36_clk _00645_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _01672_ _01677_ _01570_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _02113_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__buf_6
XFILLER_93_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07611_ _02232_ _02234_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__xnor2_4
XFILLER_81_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08591_ sha256cu.m_out_digest.b_in\[13\] _02370_ _02110_ _02027_ VGND VGND VPWR VPWR
+ _00140_ sky130_fd_sc_hd__o22a_1
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07542_ _02127_ _02131_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__o21a_1
X_07473_ _02071_ _02100_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09212_ sha256cu.m_out_digest.e_in\[19\] _02040_ _03694_ _02068_ VGND VGND VPWR VPWR
+ _00242_ sky130_fd_sc_hd__a211o_1
XFILLER_50_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09143_ _03622_ _03626_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__and2_1
XFILLER_147_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09074_ sha256cu.m_out_digest.h_in\[15\] sha256cu.m_out_digest.d_in\[15\] VGND VGND
+ VPWR VPWR _03561_ sky130_fd_sc_hd__or2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08025_ sha256cu.m_out_digest.b_in\[17\] _02162_ _02637_ VGND VGND VPWR VPWR _02638_
+ sky130_fd_sc_hd__o21ai_1
Xpassword_cracker_268 VGND VGND VPWR VPWR password_cracker_268/HI password_count[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_150_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xpassword_cracker_279 VGND VGND VPWR VPWR password_cracker_279/HI password_count[19]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09976_ sha256cu.msg_scheduler.mreg_0\[24\] _04221_ _04222_ _04211_ VGND VGND VPWR
+ VPWR _00484_ sky130_fd_sc_hd__o211a_1
XFILLER_89_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08927_ _02002_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__or2_1
X_08858_ _02230_ _03324_ _03323_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07809_ _02378_ _02389_ _02427_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__o21ba_1
X_08789_ _03263_ _03285_ _02439_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__o21ai_1
X_10820_ sha256cu.m_pad_pars.m_size\[3\] _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__or2_1
XFILLER_26_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10751_ sha256cu.msg_scheduler.mreg_11\[5\] _04659_ _04664_ _04662_ VGND VGND VPWR
+ VPWR _00817_ sky130_fd_sc_hd__o211a_1
XFILLER_41_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13470_ _06745_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_1
X_10682_ sha256cu.msg_scheduler.mreg_10\[7\] _04620_ _04625_ _04623_ VGND VGND VPWR
+ VPWR _00787_ sky130_fd_sc_hd__o211a_1
XFILLER_71_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12421_ sha256cu.m_pad_pars.block_512\[4\]\[2\] _06178_ VGND VGND VPWR VPWR _06181_
+ sky130_fd_sc_hd__and2_1
XFILLER_9_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12352_ _06145_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
X_12283_ _06085_ _06086_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__nor2_2
XFILLER_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11303_ _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__clkbuf_4
X_14022_ clknet_leaf_56_clk _00568_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11234_ _04753_ _04794_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__nor2_1
XFILLER_5_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11165_ sha256cu.m_pad_pars.block_512\[22\]\[1\] _05013_ _04977_ sha256cu.m_pad_pars.block_512\[46\]\[1\]
+ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__a221o_1
X_10116_ sha256cu.msg_scheduler.mreg_2\[20\] _04301_ _04302_ _04291_ VGND VGND VPWR
+ VPWR _00544_ sky130_fd_sc_hd__o211a_1
XFILLER_110_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11096_ _04771_ _04787_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__nor2_1
X_10047_ _01972_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__buf_2
X_14924_ clknet_leaf_10_clk _01438_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14855_ clknet_leaf_11_clk _01369_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[54\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13806_ clknet_leaf_48_clk _00352_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11998_ _05792_ _05795_ _05813_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__a21oi_1
X_14786_ clknet_leaf_107_clk _01300_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13737_ clknet_leaf_70_clk _00283_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10949_ _04815_ _04794_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_70_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_71_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13668_ clknet_leaf_87_clk _00214_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13599_ clknet_leaf_69_clk _00145_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12619_ sha256cu.m_pad_pars.block_512\[15\]\[6\] _06280_ VGND VGND VPWR VPWR _06287_
+ sky130_fd_sc_hd__and2_1
XFILLER_129_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09830_ sha256cu.msg_scheduler.mreg_13\[3\] _04134_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__or2_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09761_ sha256cu.msg_scheduler.mreg_14\[6\] _04093_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__or2_1
XFILLER_86_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _01657_ _01658_ _01659_ _01661_ _01617_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__o311a_1
XFILLER_132_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08712_ sha256cu.iter_processing.w\[1\] _02045_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__or2_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09692_ sha256cu.iter_processing.w\[8\] _04054_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__or2_1
XFILLER_67_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08643_ sha256cu.m_out_digest.c_in\[23\] _03184_ _03182_ sha256cu.m_out_digest.b_in\[23\]
+ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__a22o_1
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08574_ _03142_ _03145_ _03172_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__a21oi_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ sha256cu.m_out_digest.b_in\[4\] sha256cu.m_out_digest.a_in\[4\] VGND VGND
+ VPWR VPWR _02151_ sky130_fd_sc_hd__or2_1
XFILLER_41_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07456_ sha256cu.m_out_digest.a_in\[15\] VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07387_ _01564_ _02016_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__nand2_4
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09126_ _03502_ _03554_ _03609_ _03611_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__o31a_1
XFILLER_135_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09057_ _03540_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__xor2_1
XFILLER_108_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08008_ _02585_ _02545_ _02583_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__nor3b_2
XFILLER_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09959_ sha256cu.msg_scheduler.mreg_1\[17\] _04202_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__or2_1
XFILLER_89_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12970_ sha256cu.m_pad_pars.block_512\[36\]\[2\] _06471_ VGND VGND VPWR VPWR _06474_
+ sky130_fd_sc_hd__and2_1
XANTENNA_401 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _05738_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__and2_1
XFILLER_45_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _05642_ _05646_ _05643_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__a21boi_1
XFILLER_72_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14640_ clknet_leaf_2_clk _01154_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_412 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ sha256cu.msg_scheduler.mreg_12\[28\] _04692_ VGND VGND VPWR VPWR _04694_
+ sky130_fd_sc_hd__or2_1
X_14571_ clknet_leaf_21_clk _01085_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
X_11783_ sha256cu.msg_scheduler.mreg_14\[25\] sha256cu.msg_scheduler.mreg_14\[18\]
+ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13522_ clknet_leaf_124_clk _00072_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[63\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10734_ sha256cu.msg_scheduler.mreg_11\[30\] _04653_ VGND VGND VPWR VPWR _04655_
+ sky130_fd_sc_hd__or2_1
XFILLER_41_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10665_ sha256cu.msg_scheduler.mreg_11\[0\] _04614_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__or2_1
X_13453_ sha256cu.K\[7\] _06726_ _06727_ _06735_ _05040_ VGND VGND VPWR VPWR _01448_
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12404_ sha256cu.m_pad_pars.block_512\[3\]\[2\] _06169_ VGND VGND VPWR VPWR _06172_
+ sky130_fd_sc_hd__and2_1
X_13384_ _01923_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__buf_2
X_10596_ sha256cu.msg_scheduler.mreg_9\[2\] _04567_ _04576_ _04570_ VGND VGND VPWR
+ VPWR _00750_ sky130_fd_sc_hd__o211a_1
X_12335_ _06134_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12266_ _06042_ _06043_ _06040_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__a21oi_1
X_14005_ clknet_leaf_41_clk _00551_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_12197_ _06003_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__and2b_1
X_11217_ sha256cu.data_in_padd\[13\] _04840_ _05067_ _05070_ _05040_ VGND VGND VPWR
+ VPWR _00876_ sky130_fd_sc_hd__o221a_1
XFILLER_150_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11148_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__inv_2
XFILLER_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput170 hash[252] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xinput181 hash[31] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_2
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11079_ sha256cu.m_pad_pars.add_out3\[5\] sha256cu.m_pad_pars.add_out3\[4\] _04730_
+ _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__or4_1
XFILLER_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput192 hash[41] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14907_ clknet_leaf_125_clk _01421_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14838_ clknet_leaf_10_clk _01352_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07310_ sha256cu.byte_stop _01952_ _01953_ sha256cu.m_pad_pars.add_512_block\[1\]
+ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__or4b_1
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14769_ clknet_leaf_2_clk _01283_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08290_ _02893_ _02895_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07241_ _01653_ _01768_ _01684_ _01763_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__a31o_1
XFILLER_145_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07172_ _01694_ _01762_ _01840_ _01703_ _01584_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__o221a_1
XFILLER_20_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09813_ sha256cu.msg_scheduler.mreg_14\[28\] _04120_ VGND VGND VPWR VPWR _04127_
+ sky130_fd_sc_hd__or2_1
XFILLER_86_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09744_ sha256cu.msg_scheduler.mreg_14\[30\] _04086_ _04087_ _04077_ VGND VGND VPWR
+ VPWR _00381_ sky130_fd_sc_hd__o211a_1
X_06956_ _01590_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_4
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09675_ sha256cu.iter_processing.w\[1\] _04046_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__or2_1
X_06887_ _01578_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__nor2_1
XFILLER_27_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08626_ sha256cu.m_out_digest.c_in\[10\] _03179_ _03178_ sha256cu.m_out_digest.b_in\[10\]
+ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__a22o_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
X_08557_ sha256cu.m_out_digest.e_in\[10\] sha256cu.m_out_digest.e_in\[5\] VGND VGND
+ VPWR VPWR _03156_ sky130_fd_sc_hd__xnor2_4
XFILLER_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07508_ _02132_ _02134_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__xnor2_1
X_08488_ sha256cu.m_out_digest.g_in\[29\] sha256cu.m_out_digest.f_in\[29\] sha256cu.m_out_digest.e_in\[29\]
+ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__mux2_2
X_07439_ _02002_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__buf_6
X_10450_ sha256cu.msg_scheduler.mreg_8\[4\] _04481_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__or2_1
XFILLER_6_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09109_ _03593_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__nor2_1
X_10381_ sha256cu.msg_scheduler.mreg_7\[6\] _04441_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__or2_1
XFILLER_123_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12120_ _05929_ _05930_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__nor2_1
XFILLER_2_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12051_ _05862_ _05863_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11002_ sha256cu.m_pad_pars.block_512\[3\]\[3\] _04765_ _04774_ sha256cu.m_pad_pars.block_512\[7\]\[3\]
+ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a22o_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12953_ sha256cu.m_pad_pars.block_512\[35\]\[2\] _06462_ VGND VGND VPWR VPWR _06465_
+ sky130_fd_sc_hd__and2_1
X_11904_ _05695_ _05700_ _05723_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__and3_1
XFILLER_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_242 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_231 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14623_ clknet_leaf_97_clk _01137_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[25\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12884_ sha256cu.m_pad_pars.block_512\[31\]\[2\] _06425_ VGND VGND VPWR VPWR _06428_
+ sky130_fd_sc_hd__and2_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _05656_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__or2_1
XANTENNA_264 net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_253 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_275 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11766_ sha256cu.iter_processing.w\[7\] _05430_ _05591_ _05335_ VGND VGND VPWR VPWR
+ _00905_ sky130_fd_sc_hd__o211a_1
X_14554_ clknet_leaf_118_clk _01068_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10717_ sha256cu.msg_scheduler.mreg_11\[23\] _04640_ VGND VGND VPWR VPWR _04645_
+ sky130_fd_sc_hd__or2_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ clknet_leaf_4_clk _00999_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13505_ _06767_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_1
X_11697_ _05524_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__and2b_1
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13436_ sha256cu.K\[2\] _06714_ _06719_ _00058_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__a22o_1
X_10648_ sha256cu.msg_scheduler.mreg_10\[25\] _04601_ VGND VGND VPWR VPWR _04606_
+ sky130_fd_sc_hd__or2_1
X_10579_ sha256cu.msg_scheduler.mreg_8\[27\] _04554_ _04566_ _04557_ VGND VGND VPWR
+ VPWR _00743_ sky130_fd_sc_hd__o211a_1
XFILLER_61_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13367_ _06684_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_1
X_12318_ sha256cu.msg_scheduler.mreg_1\[17\] _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13298_ _06648_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12249_ _05963_ _05966_ _06027_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__a211o_1
XFILLER_123_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07790_ sha256cu.K\[10\] _02397_ _02408_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__a21boi_2
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06810_ net130 net133 net132 net136 VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__or4_1
XFILLER_83_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09460_ _03932_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__nor2_1
XFILLER_92_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08411_ _02967_ _02965_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_16_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
X_09391_ sha256cu.m_out_digest.e_in\[25\] _02439_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__or2_1
XFILLER_24_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08342_ sha256cu.iter_processing.w\[24\] _02904_ _02946_ VGND VGND VPWR VPWR _02947_
+ sky130_fd_sc_hd__a21oi_1
X_08273_ _02623_ _02626_ _02763_ _02878_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__a211o_1
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07224_ _01650_ _01745_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__or3_1
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07155_ _00456_ _01610_ _01773_ _01823_ _01825_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__a32o_1
XFILLER_133_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07086_ _01721_ _01701_ _01621_ _01616_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__a211o_1
XFILLER_121_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07988_ _02272_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__xnor2_2
XFILLER_86_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09727_ sha256cu.iter_processing.w\[23\] _04067_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__or2_1
X_06939_ _01621_ _01624_ _01628_ _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__o31a_1
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09658_ sha256cu.m_out_digest.h_in\[22\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[22\]
+ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__o22a_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09589_ sha256cu.m_out_digest.f_in\[28\] _04027_ _04030_ sha256cu.m_out_digest.e_in\[28\]
+ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__o22a_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08609_ sha256cu.m_out_digest.b_in\[27\] _03177_ _03176_ sha256cu.m_out_digest.a_in\[27\]
+ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__o22a_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11620_ sha256cu.msg_scheduler.mreg_1\[8\] sha256cu.msg_scheduler.mreg_1\[4\] VGND
+ VGND VPWR VPWR _05452_ sky130_fd_sc_hd__xnor2_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _05010_ _05248_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__nor2_1
X_10502_ sha256cu.msg_scheduler.mreg_7\[26\] _04513_ _04522_ _04516_ VGND VGND VPWR
+ VPWR _00710_ sky130_fd_sc_hd__o211a_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14270_ clknet_leaf_19_clk _00816_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_11\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11482_ sha256cu.data_in_padd\[24\] _01980_ _01987_ _05324_ VGND VGND VPWR VPWR _00887_
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10433_ sha256cu.msg_scheduler.mreg_6\[28\] _04474_ _04483_ _04477_ VGND VGND VPWR
+ VPWR _00680_ sky130_fd_sc_hd__o211a_1
X_13221_ _06607_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10364_ sha256cu.msg_scheduler.mreg_6\[31\] _04441_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__or2_1
X_13152_ _06570_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12103_ _05442_ _05913_ _05914_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__a21o_1
XFILLER_3_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10295_ sha256cu.msg_scheduler.mreg_5\[1\] _04393_ _04404_ _04397_ VGND VGND VPWR
+ VPWR _00621_ sky130_fd_sc_hd__o211a_1
XFILLER_97_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13083_ _06533_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__clkbuf_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12034_ sha256cu.msg_scheduler.mreg_1\[22\] sha256cu.msg_scheduler.mreg_1\[5\] VGND
+ VGND VPWR VPWR _05848_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13985_ clknet_leaf_57_clk _00531_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12936_ sha256cu.m_pad_pars.block_512\[34\]\[2\] _06453_ VGND VGND VPWR VPWR _06456_
+ sky130_fd_sc_hd__and2_1
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12867_ sha256cu.m_pad_pars.block_512\[30\]\[2\] _06416_ VGND VGND VPWR VPWR _06419_
+ sky130_fd_sc_hd__and2_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _05620_ _05635_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__and2_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14606_ clknet_leaf_110_clk _01120_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ clknet_leaf_12_clk _01051_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12798_ _06382_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11749_ _05572_ _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__xor2_1
X_14468_ clknet_leaf_100_clk _00982_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14399_ clknet_leaf_75_clk _00913_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[15\]
+ sky130_fd_sc_hd__dfxtp_4
X_13419_ sha256cu.m_pad_pars.block_512\[62\]\[6\] _01928_ VGND VGND VPWR VPWR _06711_
+ sky130_fd_sc_hd__and2_1
XFILLER_6_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08960_ _03438_ _03439_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nand2_1
XFILLER_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
X_08891_ _03382_ _03384_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__xnor2_1
X_07911_ _02128_ sha256cu.m_out_digest.a_in\[4\] VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__xnor2_1
X_07842_ _02422_ _02424_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__nor2_1
XFILLER_69_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07773_ _02390_ _02392_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__xnor2_1
X_09512_ _03951_ _03978_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__and2_1
XFILLER_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09443_ _03916_ _03917_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09374_ sha256cu.iter_processing.w\[25\] _02939_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__or2_1
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08325_ sha256cu.m_out_digest.e_in\[18\] sha256cu.m_out_digest.e_in\[4\] VGND VGND
+ VPWR VPWR _02930_ sky130_fd_sc_hd__xnor2_4
XFILLER_138_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08256_ _02815_ _02812_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__and2b_1
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08187_ sha256cu.K\[21\] _02795_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__or2_1
X_07207_ _00457_ _01865_ _01867_ _01870_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a31o_1
X_07138_ _01811_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07069_ _00454_ _01600_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__or2_1
X_10080_ _04281_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__clkbuf_2
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13770_ clknet_leaf_82_clk _00316_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10982_ sha256cu.m_pad_pars.block_512\[43\]\[1\] _04804_ _04847_ VGND VGND VPWR VPWR
+ _04848_ sky130_fd_sc_hd__a21o_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12721_ sha256cu.m_pad_pars.block_512\[21\]\[6\] _06334_ VGND VGND VPWR VPWR _06341_
+ sky130_fd_sc_hd__and2_1
XFILLER_71_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12652_ _06304_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__clkbuf_1
X_11603_ _05434_ _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__nand2_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12583_ _06267_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11534_ sha256cu.m_pad_pars.block_512\[52\]\[5\] _05310_ _05371_ _01920_ VGND VGND
+ VPWR VPWR _05372_ sky130_fd_sc_hd__a22o_1
X_14322_ clknet_leaf_90_clk _00016_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__dfxtp_1
X_14253_ clknet_leaf_25_clk _00799_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11465_ _01952_ _04761_ _05307_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__o21ai_1
X_10416_ sha256cu.msg_scheduler.mreg_6\[21\] _04461_ _04473_ _04464_ VGND VGND VPWR
+ VPWR _00673_ sky130_fd_sc_hd__o211a_1
XFILLER_143_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13204_ _06598_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_1
X_14184_ clknet_leaf_29_clk _00730_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11396_ _01985_ _05152_ _05236_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__a31o_1
X_10347_ _04314_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__clkbuf_4
XFILLER_125_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13135_ _06561_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10278_ sha256cu.msg_scheduler.mreg_4\[26\] _04393_ _04394_ _04383_ VGND VGND VPWR
+ VPWR _00614_ sky130_fd_sc_hd__o211a_1
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _06524_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__clkbuf_1
X_12017_ sha256cu.msg_scheduler.mreg_14\[28\] _05831_ VGND VGND VPWR VPWR _05832_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_48_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13968_ clknet_leaf_54_clk _00514_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[22\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_62_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12919_ sha256cu.m_pad_pars.block_512\[33\]\[2\] _06444_ VGND VGND VPWR VPWR _06447_
+ sky130_fd_sc_hd__and2_1
X_13899_ clknet_leaf_20_clk _00445_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09090_ sha256cu.K\[14\] _03543_ _03542_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__a21o_1
X_08110_ _02710_ _02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__xor2_1
X_08041_ _02604_ _02606_ _02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__o21a_1
XFILLER_143_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09992_ sha256cu.msg_scheduler.mreg_0\[31\] _04221_ _04231_ _04224_ VGND VGND VPWR
+ VPWR _00491_ sky130_fd_sc_hd__o211a_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08943_ _03431_ _03434_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__xnor2_2
XFILLER_131_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
X_08874_ sha256cu.K\[7\] _03346_ _03345_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__a21bo_1
XFILLER_96_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07825_ sha256cu.iter_processing.w\[11\] _02414_ _02442_ VGND VGND VPWR VPWR _02443_
+ sky130_fd_sc_hd__a21o_1
XFILLER_111_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07756_ _02372_ _02373_ _02374_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__a21o_1
X_07687_ sha256cu.m_out_digest.h_in\[7\] _02275_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__nand2_1
X_09426_ _03899_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__nand2_1
XFILLER_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09357_ _03779_ _03809_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__nand2_1
XFILLER_100_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ sha256cu.K\[22\] _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08308_ _02912_ _02913_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__or2_1
X_08239_ _02818_ _02819_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__and2b_1
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11250_ _04908_ _04974_ _05101_ sha256cu.m_pad_pars.block_512\[30\]\[7\] VGND VGND
+ VPWR VPWR _05102_ sky130_fd_sc_hd__a22o_1
X_10201_ sha256cu.msg_scheduler.mreg_4\[25\] _04348_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__or2_1
XFILLER_107_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11181_ sha256cu.m_pad_pars.block_512\[50\]\[2\] _05008_ _04972_ sha256cu.m_pad_pars.block_512\[38\]\[2\]
+ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__a221o_1
X_10132_ sha256cu.msg_scheduler.mreg_2\[27\] _04301_ _04311_ _04304_ VGND VGND VPWR
+ VPWR _00551_ sky130_fd_sc_hd__o211a_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10063_ sha256cu.msg_scheduler.mreg_2\[30\] _04268_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__or2_1
XFILLER_121_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14940_ clknet_leaf_91_clk _01454_ VGND VGND VPWR VPWR sha256cu.K\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14871_ clknet_leaf_124_clk _01385_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[56\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13822_ clknet_leaf_48_clk _00368_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_63_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13753_ clknet_leaf_64_clk _00299_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10965_ _01917_ _01951_ _04771_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__or3_1
X_12704_ sha256cu.m_pad_pars.block_512\[20\]\[6\] _06325_ VGND VGND VPWR VPWR _06332_
+ sky130_fd_sc_hd__and2_1
X_13684_ clknet_leaf_65_clk _00230_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[7\]
+ sky130_fd_sc_hd__dfxtp_4
X_10896_ _01943_ _04759_ _04762_ _04698_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12635_ _06295_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12566_ _06258_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11517_ sha256cu.m_pad_pars.block_512\[24\]\[4\] _05279_ _05313_ sha256cu.m_pad_pars.block_512\[4\]\[4\]
+ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__a22o_1
X_14305_ clknet_leaf_95_clk _00029_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12497_ sha256cu.m_pad_pars.block_512\[8\]\[6\] _06214_ VGND VGND VPWR VPWR _06221_
+ sky130_fd_sc_hd__and2_1
X_14236_ clknet_leaf_19_clk _00782_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11448_ _04701_ _05154_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__nor2_1
XFILLER_152_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14167_ clknet_leaf_34_clk _00713_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11379_ sha256cu.m_pad_pars.block_512\[61\]\[6\] _05162_ _05163_ sha256cu.m_pad_pars.block_512\[57\]\[6\]
+ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__a22o_1
XFILLER_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _06552_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__clkbuf_1
X_14098_ clknet_leaf_33_clk _00644_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _06515_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08590_ sha256cu.m_out_digest.b_in\[12\] _03031_ _02114_ _02382_ VGND VGND VPWR VPWR
+ _00139_ sky130_fd_sc_hd__a22o_1
XFILLER_93_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07610_ _02233_ sha256cu.m_out_digest.a_in\[8\] VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__xnor2_2
XFILLER_81_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07541_ sha256cu.m_out_digest.h_in\[3\] _02130_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__nand2_1
XFILLER_53_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07472_ _02096_ _02099_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__xor2_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09211_ _03691_ _03692_ _03693_ _02732_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__a211oi_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09142_ _03622_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__nor2_1
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09073_ _03548_ _03549_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__nand2_1
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08024_ sha256cu.m_out_digest.b_in\[17\] _02162_ sha256cu.m_out_digest.c_in\[17\]
+ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__a21o_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpassword_cracker_269 VGND VGND VPWR VPWR password_cracker_269/HI password_count[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09975_ sha256cu.msg_scheduler.mreg_1\[24\] _04215_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__or2_1
XFILLER_104_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08926_ sha256cu.m_out_digest.e_in\[9\] _02037_ _02017_ _03418_ VGND VGND VPWR VPWR
+ _03419_ sky130_fd_sc_hd__a22o_1
X_08857_ _02270_ _03351_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__xor2_1
XFILLER_84_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07808_ _02386_ _02388_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__nor2_1
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08788_ _03263_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__and2_1
XFILLER_72_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07739_ _02357_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__xor2_1
XFILLER_60_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10750_ sha256cu.msg_scheduler.mreg_12\[5\] _04653_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__or2_1
XFILLER_41_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10681_ sha256cu.msg_scheduler.mreg_11\[7\] _04614_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__or2_1
X_09409_ _03883_ _03884_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__and2_1
XFILLER_41_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12420_ _06180_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12351_ sha256cu.m_pad_pars.block_512\[0\]\[0\] _06144_ VGND VGND VPWR VPWR _06145_
+ sky130_fd_sc_hd__and2_1
XFILLER_153_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12282_ _06083_ _06084_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__and2_1
X_11302_ _01941_ _01953_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__or2_1
X_14021_ clknet_leaf_57_clk _00567_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11233_ _04917_ _04954_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__o21a_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11164_ sha256cu.m_pad_pars.block_512\[18\]\[1\] _05014_ _05009_ sha256cu.m_pad_pars.block_512\[30\]\[1\]
+ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__a22o_1
XFILLER_49_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10115_ sha256cu.msg_scheduler.mreg_3\[20\] _04295_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__or2_1
X_11095_ _01953_ _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__or2_4
X_10046_ sha256cu.msg_scheduler.mreg_2\[23\] _04254_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__or2_1
X_14923_ clknet_leaf_9_clk _01437_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14854_ clknet_leaf_102_clk _01368_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13805_ clknet_leaf_49_clk _00351_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11997_ _05811_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__and2b_1
X_14785_ clknet_leaf_108_clk _01299_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13736_ clknet_leaf_83_clk _00282_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10948_ _04748_ _01940_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__or2_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13667_ clknet_leaf_87_clk _00213_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10879_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_129_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13598_ clknet_leaf_69_clk _00144_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12618_ _06286_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12549_ _06248_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _01479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14219_ clknet_leaf_30_clk _00765_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09760_ sha256cu.msg_scheduler.mreg_13\[5\] _04086_ _04096_ _04090_ VGND VGND VPWR
+ VPWR _00388_ sky130_fd_sc_hd__o211a_1
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _01660_ _01634_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__nand2_2
XFILLER_100_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09691_ sha256cu.msg_scheduler.mreg_14\[7\] _04045_ _04057_ _04050_ VGND VGND VPWR
+ VPWR _00358_ sky130_fd_sc_hd__o211a_1
X_08711_ sha256cu.iter_processing.w\[1\] _02045_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__nand2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08642_ sha256cu.m_out_digest.c_in\[22\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[22\]
+ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__o22a_1
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08573_ _03148_ _03171_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__xnor2_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07524_ sha256cu.iter_processing.w\[3\] _02122_ _02121_ VGND VGND VPWR VPWR _02150_
+ sky130_fd_sc_hd__a21o_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07455_ sha256cu.m_out_digest.a_in\[24\] VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__buf_4
XFILLER_50_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07386_ _02005_ _02015_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__or2_2
XFILLER_41_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09125_ _03553_ _03555_ _03581_ _03610_ _03580_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__a311oi_1
X_09056_ sha256cu.K\[14\] _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__xnor2_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08007_ _02619_ _02620_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__or2_1
XFILLER_104_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09958_ sha256cu.msg_scheduler.mreg_0\[16\] _04208_ _04212_ _04211_ VGND VGND VPWR
+ VPWR _00476_ sky130_fd_sc_hd__o211a_1
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08909_ _03399_ _03400_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__nand2_1
XFILLER_106_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09889_ _04116_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__buf_6
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11920_ _05736_ _05737_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__nand2_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _05670_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__xor2_1
XANTENNA_413 net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_402 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11782_ _05605_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__and2_1
X_10802_ sha256cu.msg_scheduler.mreg_11\[27\] _04685_ _04693_ _04688_ VGND VGND VPWR
+ VPWR _00839_ sky130_fd_sc_hd__o211a_1
XFILLER_82_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14570_ clknet_leaf_16_clk _01084_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ sha256cu.msg_scheduler.mreg_10\[29\] _04646_ _04654_ _04649_ VGND VGND VPWR
+ VPWR _00809_ sky130_fd_sc_hd__o211a_1
XFILLER_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13521_ clknet_leaf_79_clk _00071_ VGND VGND VPWR VPWR sha256cu.iter_processing.rst
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10664_ sha256cu.msg_scheduler.mreg_9\[31\] _04607_ _04615_ _04610_ VGND VGND VPWR
+ VPWR _00779_ sky130_fd_sc_hd__o211a_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13452_ _04188_ _00065_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__and2b_1
X_10595_ sha256cu.msg_scheduler.mreg_10\[2\] _04574_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__or2_1
X_12403_ _06171_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__clkbuf_1
X_13383_ _06692_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12334_ _06132_ _01983_ _06133_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__and3b_1
XFILLER_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14004_ clknet_leaf_40_clk _00550_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12265_ _06068_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nand2_1
X_12196_ _05975_ _05988_ _06002_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__a21o_1
X_11216_ sha256cu.m_pad_pars.block_512\[22\]\[5\] _05013_ _05069_ _01970_ VGND VGND
+ VPWR VPWR _05070_ sky130_fd_sc_hd__a211o_1
XFILLER_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11147_ _01952_ _05004_ _05005_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__o21bai_2
XFILLER_1_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput171 hash[253] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
X_11078_ _04937_ _04778_ _04780_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__a21bo_1
Xinput160 hash[243] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
X_10029_ sha256cu.msg_scheduler.mreg_1\[15\] _04247_ _04252_ _04250_ VGND VGND VPWR
+ VPWR _00507_ sky130_fd_sc_hd__o211a_1
Xinput182 hash[32] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
Xinput193 hash[42] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14906_ clknet_leaf_125_clk _01420_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14837_ clknet_leaf_4_clk _01351_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14768_ clknet_leaf_1_clk _01282_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13719_ clknet_leaf_65_clk _00265_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14699_ clknet_leaf_7_clk _01213_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07240_ _01724_ _01897_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__nand2_1
X_07171_ _01830_ _01658_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__nor2_1
XFILLER_117_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09812_ _04044_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__buf_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09743_ sha256cu.iter_processing.w\[30\] _04080_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__or2_1
X_06955_ _01636_ _01638_ _01641_ _01643_ _01644_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__o221a_1
X_09674_ sha256cu.msg_scheduler.mreg_14\[0\] _04045_ _04047_ _03366_ VGND VGND VPWR
+ VPWR _00351_ sky130_fd_sc_hd__o211a_1
XFILLER_55_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06886_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__buf_4
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08625_ sha256cu.m_out_digest.c_in\[9\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[9\]
+ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__o22a_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08556_ sha256cu.iter_processing.w\[30\] _03127_ _03154_ VGND VGND VPWR VPWR _03155_
+ sky130_fd_sc_hd__a21oi_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07507_ _02082_ _02087_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__o21a_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08487_ sha256cu.m_out_digest.b_in\[29\] _02272_ _03087_ VGND VGND VPWR VPWR _03088_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07438_ _02035_ _02063_ _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__o21a_1
XFILLER_10_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07369_ sha256cu.counter_iteration\[5\] sha256cu.counter_iteration\[4\] sha256cu.counter_iteration\[6\]
+ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__or3b_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09108_ sha256cu.iter_processing.w\[16\] _02595_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__and2_1
XFILLER_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10380_ sha256cu.msg_scheduler.mreg_6\[5\] _04448_ _04453_ _04451_ VGND VGND VPWR
+ VPWR _00657_ sky130_fd_sc_hd__o211a_1
XFILLER_117_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09039_ _03496_ _03503_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12050_ sha256cu.data_in_padd\[19\] _05667_ _05445_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11001_ sha256cu.m_pad_pars.block_512\[27\]\[3\] _04757_ _04804_ sha256cu.m_pad_pars.block_512\[43\]\[3\]
+ _04864_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__a221o_1
XFILLER_132_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12952_ _06464_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__clkbuf_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _05720_ _05722_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__xnor2_1
XANTENNA_243 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_232 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_210 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14622_ clknet_leaf_115_clk _01136_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12883_ _06427_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__clkbuf_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _05630_ _05632_ _05628_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__a21oi_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_254 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_287 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ sha256cu.data_in_padd\[7\] _05448_ _05590_ _05463_ VGND VGND VPWR VPWR _05591_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_298 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14553_ clknet_leaf_119_clk _01067_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10716_ sha256cu.msg_scheduler.mreg_10\[22\] _04633_ _04644_ _04636_ VGND VGND VPWR
+ VPWR _00802_ sky130_fd_sc_hd__o211a_1
X_11696_ _05506_ _05502_ _05523_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__a21o_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14484_ clknet_leaf_5_clk _00998_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13504_ _01975_ _06766_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__and2_1
X_10647_ sha256cu.msg_scheduler.mreg_9\[24\] _04594_ _04605_ _04597_ VGND VGND VPWR
+ VPWR _00772_ sky130_fd_sc_hd__o211a_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13435_ _06723_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10578_ sha256cu.msg_scheduler.mreg_9\[27\] _04561_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__or2_1
X_13366_ sha256cu.m_pad_pars.block_512\[59\]\[4\] _06682_ VGND VGND VPWR VPWR _06684_
+ sky130_fd_sc_hd__and2_1
X_12317_ sha256cu.msg_scheduler.mreg_14\[18\] sha256cu.msg_scheduler.mreg_14\[16\]
+ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__xnor2_1
X_13297_ sha256cu.m_pad_pars.block_512\[55\]\[3\] _06644_ VGND VGND VPWR VPWR _06648_
+ sky130_fd_sc_hd__and2_1
XFILLER_142_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12248_ _06026_ _06046_ _06047_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__or3_1
XFILLER_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12179_ sha256cu.iter_processing.w\[24\] _05894_ _05987_ _05866_ VGND VGND VPWR VPWR
+ _00922_ sky130_fd_sc_hd__o211a_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08410_ _03011_ _03012_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__nand2_1
X_09390_ _03832_ _03840_ _03865_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08341_ _02902_ _02903_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__and2b_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08272_ _02839_ _02840_ _02874_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__or3_1
X_07223_ _01593_ _01648_ _01647_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07154_ _01601_ _01658_ _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__or3b_1
X_07085_ _01761_ _01763_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__or2_1
XFILLER_101_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07987_ _02198_ sha256cu.m_out_digest.a_in\[6\] VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09726_ sha256cu.msg_scheduler.mreg_14\[22\] _04073_ _04076_ _04077_ VGND VGND VPWR
+ VPWR _00373_ sky130_fd_sc_hd__o211a_1
X_06938_ _01571_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09657_ sha256cu.m_out_digest.h_in\[21\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[21\]
+ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__o22a_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06869_ sha256cu.iter_processing.rst VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__buf_8
XFILLER_28_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09588_ _02109_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__buf_4
XFILLER_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08608_ sha256cu.m_out_digest.b_in\[26\] _03179_ _03178_ _02161_ VGND VGND VPWR VPWR
+ _00153_ sky130_fd_sc_hd__a22o_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _03095_ _03113_ _03137_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__or3b_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11550_ _05314_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__inv_2
X_10501_ sha256cu.msg_scheduler.mreg_8\[26\] _04520_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__or2_1
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13220_ sha256cu.m_pad_pars.block_512\[50\]\[7\] _05109_ _06542_ VGND VGND VPWR VPWR
+ _06607_ sky130_fd_sc_hd__mux2_1
X_11481_ _05290_ _05301_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__or3_2
X_10432_ sha256cu.msg_scheduler.mreg_7\[28\] _04481_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__or2_1
XFILLER_152_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10363_ sha256cu.msg_scheduler.mreg_5\[30\] _04434_ _04443_ _04437_ VGND VGND VPWR
+ VPWR _00650_ sky130_fd_sc_hd__o211a_1
XFILLER_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13151_ sha256cu.m_pad_pars.block_512\[46\]\[7\] _05113_ _06542_ VGND VGND VPWR VPWR
+ _06570_ sky130_fd_sc_hd__mux2_1
X_12102_ sha256cu.data_in_padd\[21\] _05447_ _04692_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__a21o_1
X_13082_ sha256cu.m_pad_pars.block_512\[42\]\[7\] _05087_ _06442_ VGND VGND VPWR VPWR
+ _06533_ sky130_fd_sc_hd__mux2_1
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10294_ sha256cu.msg_scheduler.mreg_6\[1\] _04401_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__or2_1
X_12033_ _05845_ _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__nand2_1
XFILLER_78_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13984_ clknet_leaf_56_clk _00530_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12935_ _06455_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__clkbuf_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _06418_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__clkbuf_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ sha256cu.iter_processing.w\[9\] _05430_ _05639_ _05640_ VGND VGND VPWR VPWR
+ _00907_ sky130_fd_sc_hd__o211a_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ clknet_leaf_15_clk _01119_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ clknet_leaf_12_clk _01050_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12797_ sha256cu.m_pad_pars.block_512\[26\]\[1\] _06380_ VGND VGND VPWR VPWR _06382_
+ sky130_fd_sc_hd__and2_1
XFILLER_42_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11748_ sha256cu.msg_scheduler.mreg_1\[25\] _05573_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__xnor2_1
X_11679_ sha256cu.msg_scheduler.mreg_9\[4\] sha256cu.msg_scheduler.mreg_0\[4\] VGND
+ VGND VPWR VPWR _05508_ sky130_fd_sc_hd__or2_1
X_14467_ clknet_leaf_98_clk _00981_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14398_ clknet_leaf_47_clk _00912_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[14\]
+ sky130_fd_sc_hd__dfxtp_4
X_13418_ _06710_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_1
X_13349_ sha256cu.m_pad_pars.block_512\[58\]\[4\] _06671_ VGND VGND VPWR VPWR _06675_
+ sky130_fd_sc_hd__and2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08890_ _03348_ _03354_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__o21a_1
XFILLER_123_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07910_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__inv_2
XFILLER_68_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07841_ _02448_ _02458_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__xor2_1
X_07772_ _02342_ _02352_ _02391_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__o21ba_1
X_09511_ sha256cu.m_out_digest.e_in\[29\] _02440_ _03982_ _03983_ _01974_ VGND VGND
+ VPWR VPWR _00252_ sky130_fd_sc_hd__o221a_1
XFILLER_56_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09442_ sha256cu.K\[26\] _03880_ _03879_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__a21o_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09373_ _03848_ _03849_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__or2_1
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08324_ sha256cu.m_out_digest.h_in\[25\] _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08255_ _02856_ _02861_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__xnor2_1
X_08186_ _02792_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__xnor2_1
X_07206_ _01745_ _01831_ _01869_ _01663_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__o211a_1
XFILLER_119_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07137_ _01807_ _01810_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__or2_1
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07068_ _01747_ _01748_ _01644_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09709_ sha256cu.iter_processing.w\[15\] _04067_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__or2_1
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10981_ sha256cu.m_pad_pars.block_512\[59\]\[1\] _04829_ _04822_ sha256cu.m_pad_pars.block_512\[47\]\[1\]
+ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__a22o_1
XFILLER_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12720_ _06340_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12651_ sha256cu.m_pad_pars.block_512\[17\]\[5\] _06298_ VGND VGND VPWR VPWR _06304_
+ sky130_fd_sc_hd__and2_1
XFILLER_31_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11602_ sha256cu.msg_scheduler.mreg_9\[0\] sha256cu.msg_scheduler.mreg_0\[0\] VGND
+ VGND VPWR VPWR _05435_ sky130_fd_sc_hd__or2_1
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12582_ sha256cu.m_pad_pars.block_512\[13\]\[5\] _06261_ VGND VGND VPWR VPWR _06267_
+ sky130_fd_sc_hd__and2_1
XFILLER_11_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11533_ sha256cu.m_pad_pars.block_512\[60\]\[5\] _01998_ _05280_ sha256cu.m_pad_pars.block_512\[56\]\[5\]
+ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__a22o_1
X_14321_ clknet_leaf_89_clk _00015_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__dfxtp_1
X_14252_ clknet_leaf_26_clk _00798_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11464_ _04703_ _04824_ _05154_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__or3_1
X_10415_ sha256cu.msg_scheduler.mreg_7\[21\] _04468_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__or2_1
XFILLER_109_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13203_ sha256cu.m_pad_pars.block_512\[49\]\[7\] _05270_ _06542_ VGND VGND VPWR VPWR
+ _06598_ sky130_fd_sc_hd__mux2_1
X_14183_ clknet_leaf_29_clk _00729_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11395_ _05127_ _05152_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__and3_1
X_10346_ sha256cu.msg_scheduler.mreg_5\[23\] _04421_ _04433_ _04424_ VGND VGND VPWR
+ VPWR _00643_ sky130_fd_sc_hd__o211a_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13134_ sha256cu.m_pad_pars.block_512\[45\]\[7\] _05256_ _06542_ VGND VGND VPWR VPWR
+ _06561_ sky130_fd_sc_hd__mux2_1
X_10277_ sha256cu.msg_scheduler.mreg_5\[26\] _04387_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__or2_1
XFILLER_105_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ sha256cu.m_pad_pars.block_512\[41\]\[7\] _05232_ _06442_ VGND VGND VPWR VPWR
+ _06524_ sky130_fd_sc_hd__mux2_1
X_12016_ sha256cu.msg_scheduler.mreg_14\[5\] sha256cu.msg_scheduler.mreg_14\[3\] VGND
+ VGND VPWR VPWR _05831_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13967_ clknet_leaf_55_clk _00513_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[21\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12918_ _06446_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__clkbuf_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13898_ clknet_leaf_22_clk _00444_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12849_ _06409_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__clkbuf_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14519_ clknet_leaf_122_clk _01033_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08040_ _02597_ _02607_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__or2_1
XFILLER_127_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09991_ sha256cu.msg_scheduler.mreg_1\[31\] _04228_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__or2_1
XFILLER_115_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08942_ _03432_ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__nand2_1
XFILLER_131_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08873_ _03342_ _03358_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__nand2_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07824_ _02412_ _02413_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__and2b_1
XFILLER_96_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07755_ _02372_ _02373_ _02374_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__and3_1
X_07686_ _02303_ _02307_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__xnor2_2
X_09425_ sha256cu.m_out_digest.h_in\[27\] sha256cu.m_out_digest.d_in\[27\] VGND VGND
+ VPWR VPWR _03900_ sky130_fd_sc_hd__or2_1
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09356_ _03832_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__nand2_1
XFILLER_40_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09287_ _03765_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__nor2_1
X_08307_ _02862_ _02864_ _02866_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__o21ba_1
X_08238_ _02026_ _02070_ _02845_ _01984_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__a22o_1
X_10200_ sha256cu.msg_scheduler.mreg_3\[24\] _04341_ _04350_ _04344_ VGND VGND VPWR
+ VPWR _00580_ sky130_fd_sc_hd__o211a_1
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08169_ _02775_ _02777_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11180_ sha256cu.m_pad_pars.block_512\[34\]\[2\] _04996_ _04981_ sha256cu.m_pad_pars.block_512\[54\]\[2\]
+ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__a22o_1
X_10131_ sha256cu.msg_scheduler.mreg_3\[27\] _04308_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__or2_1
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10062_ sha256cu.msg_scheduler.mreg_1\[29\] _04260_ _04271_ _04264_ VGND VGND VPWR
+ VPWR _00521_ sky130_fd_sc_hd__o211a_1
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14870_ clknet_leaf_123_clk _01384_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[55\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13821_ clknet_leaf_48_clk _00367_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_75_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13752_ clknet_leaf_65_clk _00298_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10964_ _04756_ _04764_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__and3_2
X_12703_ _06331_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__clkbuf_1
X_13683_ clknet_leaf_65_clk _00229_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10895_ _01943_ _04761_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__nor2_1
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12634_ sha256cu.m_pad_pars.block_512\[16\]\[5\] _06289_ VGND VGND VPWR VPWR _06295_
+ sky130_fd_sc_hd__and2_1
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12565_ sha256cu.m_pad_pars.block_512\[12\]\[5\] _06252_ VGND VGND VPWR VPWR _06258_
+ sky130_fd_sc_hd__and2_1
X_11516_ sha256cu.data_in_padd\[27\] _01980_ _01987_ _05355_ VGND VGND VPWR VPWR _00890_
+ sky130_fd_sc_hd__a22o_1
X_14304_ clknet_leaf_90_clk _00028_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12496_ _06220_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__clkbuf_1
X_14235_ clknet_leaf_19_clk _00781_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11447_ sha256cu.m_pad_pars.block_512\[24\]\[0\] _05279_ _05281_ _01921_ _05289_
+ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__a221o_1
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14166_ clknet_leaf_34_clk _00712_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11378_ sha256cu.m_pad_pars.block_512\[1\]\[6\] _05135_ _05138_ sha256cu.m_pad_pars.block_512\[17\]\[6\]
+ _05222_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__a221o_1
X_10329_ sha256cu.msg_scheduler.mreg_5\[15\] _04421_ _04423_ _04424_ VGND VGND VPWR
+ VPWR _00635_ sky130_fd_sc_hd__o211a_1
XFILLER_124_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ sha256cu.m_pad_pars.block_512\[44\]\[7\] _05390_ _06542_ VGND VGND VPWR VPWR
+ _06552_ sky130_fd_sc_hd__mux2_1
X_14097_ clknet_leaf_33_clk _00643_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ sha256cu.m_pad_pars.block_512\[40\]\[7\] _05400_ _06442_ VGND VGND VPWR VPWR
+ _06515_ sky130_fd_sc_hd__mux2_1
XFILLER_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07540_ _02160_ _02165_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07471_ _02042_ _02097_ _02098_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09210_ _03691_ _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__nor2_1
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09141_ sha256cu.K\[17\] _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__xnor2_1
X_09072_ _02923_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__clkbuf_4
X_08023_ sha256cu.iter_processing.w\[16\] _02596_ _02635_ VGND VGND VPWR VPWR _02636_
+ sky130_fd_sc_hd__a21o_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09974_ _04166_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__clkbuf_4
XFILLER_103_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08925_ _03415_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08856_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nand2_1
XFILLER_112_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07807_ _02415_ _02425_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__xor2_2
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08787_ _03282_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__xor2_2
XFILLER_85_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07738_ _02293_ _02315_ _02358_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07669_ _02290_ _02291_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10680_ sha256cu.msg_scheduler.mreg_10\[6\] _04620_ _04624_ _04623_ VGND VGND VPWR
+ VPWR _00786_ sky130_fd_sc_hd__o211a_1
X_09408_ _03848_ _03856_ _03882_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__or3_1
XFILLER_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09339_ _02851_ _03786_ _03787_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__a21boi_1
XFILLER_153_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12350_ _01986_ _05264_ _04787_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__or3_2
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12281_ _06083_ _06084_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__nor2_1
X_11301_ sha256cu.m_pad_pars.add_out1\[3\] sha256cu.m_pad_pars.add_out1\[2\] VGND
+ VGND VPWR VPWR _05152_ sky130_fd_sc_hd__nor2b_2
X_14020_ clknet_leaf_56_clk _00566_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11232_ _04698_ _04970_ sha256cu.m_pad_pars.block_512\[38\]\[7\] VGND VGND VPWR VPWR
+ _05084_ sky130_fd_sc_hd__a21o_1
X_11163_ sha256cu.m_pad_pars.block_512\[10\]\[1\] _04963_ _04972_ sha256cu.m_pad_pars.block_512\[38\]\[1\]
+ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__a221o_1
X_10114_ _04166_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__buf_2
XFILLER_122_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11094_ sha256cu.m_pad_pars.add_512_block\[1\] _01939_ VGND VGND VPWR VPWR _04953_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10045_ sha256cu.msg_scheduler.mreg_1\[22\] _04260_ _04261_ _04250_ VGND VGND VPWR
+ VPWR _00514_ sky130_fd_sc_hd__o211a_1
X_14922_ clknet_leaf_9_clk _01436_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14853_ clknet_leaf_99_clk _01367_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13804_ clknet_leaf_70_clk _00350_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11996_ _05783_ _05788_ _05810_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__a21o_1
X_14784_ clknet_leaf_106_clk _01298_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13735_ clknet_leaf_83_clk _00281_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10947_ _04735_ sha256cu.m_pad_pars.add_out3\[4\] VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__or2_1
XFILLER_71_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13666_ clknet_leaf_87_clk _00212_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_12617_ sha256cu.m_pad_pars.block_512\[15\]\[5\] _06280_ VGND VGND VPWR VPWR _06286_
+ sky130_fd_sc_hd__and2_1
X_10878_ _04703_ _04744_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_129_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13597_ clknet_leaf_69_clk _00143_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12548_ sha256cu.m_pad_pars.block_512\[11\]\[6\] _06241_ VGND VGND VPWR VPWR _06248_
+ sky130_fd_sc_hd__and2_1
XFILLER_117_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12479_ _06211_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 _01479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14218_ clknet_leaf_30_clk _00764_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14149_ clknet_leaf_33_clk _00695_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _01586_ _01588_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__nor2_1
X_09690_ sha256cu.iter_processing.w\[7\] _04054_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__or2_1
X_08710_ sha256cu.K\[1\] VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__inv_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08641_ sha256cu.m_out_digest.c_in\[21\] _03185_ _03183_ sha256cu.m_out_digest.b_in\[21\]
+ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__o22a_1
XFILLER_39_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08572_ _03151_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__xnor2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07523_ sha256cu.m_out_digest.a_in\[3\] _02070_ _02114_ _02149_ VGND VGND VPWR VPWR
+ _00098_ sky130_fd_sc_hd__a22o_1
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07454_ _02081_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__inv_2
XFILLER_50_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07385_ sha256cu.iter_processing.temp_case sha256cu.iter_processing.padding_done
+ sha256cu.iter_processing.temp_if VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__a21oi_2
XFILLER_136_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09124_ _03551_ _03579_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__nor2_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09055_ _03541_ _03542_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__nor2_1
X_08006_ _02589_ _02590_ _02618_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__and3_1
XFILLER_151_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09957_ sha256cu.msg_scheduler.mreg_1\[16\] _04202_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__or2_1
XFILLER_89_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08908_ _03399_ _03400_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__nor2_1
X_09888_ sha256cu.msg_scheduler.mreg_13\[28\] _04160_ VGND VGND VPWR VPWR _04170_
+ sky130_fd_sc_hd__or2_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _03304_ _03305_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__a21bo_1
XFILLER_73_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ sha256cu.msg_scheduler.mreg_1\[29\] _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_403 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _05603_ _05604_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__nand2_1
X_10801_ sha256cu.msg_scheduler.mreg_12\[27\] _04692_ VGND VGND VPWR VPWR _04693_
+ sky130_fd_sc_hd__or2_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10732_ sha256cu.msg_scheduler.mreg_11\[29\] _04653_ VGND VGND VPWR VPWR _04654_
+ sky130_fd_sc_hd__or2_1
X_13520_ clknet_leaf_109_clk _00070_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dfxtp_1
XFILLER_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10663_ sha256cu.msg_scheduler.mreg_10\[31\] _04614_ VGND VGND VPWR VPWR _04615_
+ sky130_fd_sc_hd__or2_1
X_13451_ _06734_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_1
X_10594_ sha256cu.msg_scheduler.mreg_9\[1\] _04567_ _04575_ _04570_ VGND VGND VPWR
+ VPWR _00749_ sky130_fd_sc_hd__o211a_1
X_12402_ sha256cu.m_pad_pars.block_512\[3\]\[1\] _06169_ VGND VGND VPWR VPWR _06171_
+ sky130_fd_sc_hd__and2_1
X_13382_ sha256cu.m_pad_pars.block_512\[60\]\[4\] _06682_ VGND VGND VPWR VPWR _06692_
+ sky130_fd_sc_hd__and2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12333_ _01939_ _01947_ sha256cu.m_pad_pars.add_512_block\[1\] VGND VGND VPWR VPWR
+ _06133_ sky130_fd_sc_hd__a21o_1
XFILLER_142_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14003_ clknet_leaf_41_clk _00549_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12264_ _06066_ _06067_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__or2_1
XFILLER_5_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12195_ _05975_ _05988_ _06002_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__and3_1
X_11215_ sha256cu.m_pad_pars.block_512\[50\]\[5\] _05008_ _04972_ sha256cu.m_pad_pars.block_512\[38\]\[5\]
+ _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__a221o_1
XFILLER_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11146_ _04759_ _04824_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__nor2_1
XFILLER_95_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11077_ sha256cu.m_pad_pars.block_512\[15\]\[7\] VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__inv_2
X_10028_ sha256cu.msg_scheduler.mreg_2\[15\] _04241_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__or2_1
Xinput150 hash[234] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_4
Xinput172 hash[254] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
Xinput161 hash[244] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14905_ clknet_leaf_124_clk _01419_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput183 hash[33] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput194 hash[43] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14836_ clknet_leaf_1_clk _01350_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_91_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14767_ clknet_leaf_3_clk _01281_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[43\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13718_ clknet_leaf_65_clk _00264_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11979_ _05775_ _05794_ _05442_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__o21a_1
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14698_ clknet_leaf_22_clk _01212_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13649_ clknet_leaf_60_clk _00195_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07170_ _01636_ _01682_ _01729_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__o21ba_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_113_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09811_ sha256cu.msg_scheduler.mreg_13\[27\] _04112_ _04125_ _04117_ VGND VGND VPWR
+ VPWR _00410_ sky130_fd_sc_hd__o211a_1
XFILLER_101_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09742_ _04044_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__clkbuf_4
X_06954_ _01620_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09673_ sha256cu.iter_processing.w\[0\] _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__or2_1
X_06885_ sha256cu.counter_iteration\[1\] sha256cu.msg_scheduler.counter_iteration\[1\]
+ _01568_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__mux2_2
X_08624_ sha256cu.m_out_digest.c_in\[8\] _03181_ _03180_ sha256cu.m_out_digest.b_in\[8\]
+ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__o22a_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08555_ _03125_ _03126_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__and2b_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07506_ sha256cu.m_out_digest.h_in\[2\] _02086_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__nand2_1
XFILLER_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08486_ sha256cu.m_out_digest.b_in\[29\] _02272_ sha256cu.m_out_digest.c_in\[29\]
+ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__a21o_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07437_ _02035_ _02063_ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07368_ sha256cu.m_pad_pars.add_out0\[6\] _02001_ _02003_ VGND VGND VPWR VPWR _00089_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09107_ sha256cu.iter_processing.w\[16\] _02595_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__nor2_1
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_111_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_16
X_07299_ sha256cu.m_pad_pars.add_512_block\[5\] sha256cu.m_pad_pars.add_512_block\[4\]
+ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__or2_2
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09038_ _03525_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__and2b_1
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11000_ sha256cu.m_pad_pars.block_512\[51\]\[3\] _04826_ _04822_ sha256cu.m_pad_pars.block_512\[47\]\[3\]
+ _04863_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__a221o_1
XFILLER_89_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12951_ sha256cu.m_pad_pars.block_512\[35\]\[1\] _06462_ VGND VGND VPWR VPWR _06464_
+ sky130_fd_sc_hd__and2_1
XANTENNA_200 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ sha256cu.msg_scheduler.mreg_14\[30\] _05721_ VGND VGND VPWR VPWR _05722_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_73_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12882_ sha256cu.m_pad_pars.block_512\[31\]\[1\] _06425_ VGND VGND VPWR VPWR _06427_
+ sky130_fd_sc_hd__and2_1
XANTENNA_211 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_233 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11833_ _05654_ _05655_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__nand2_1
XFILLER_93_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14621_ clknet_leaf_121_clk _01135_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 sha256cu.iter_processing.w\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_255 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_266 net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _05465_ _05589_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__nor2_1
XANTENNA_299 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14552_ clknet_leaf_119_clk _01066_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10715_ sha256cu.msg_scheduler.mreg_11\[22\] _04640_ VGND VGND VPWR VPWR _04644_
+ sky130_fd_sc_hd__or2_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _05506_ _05502_ _05523_ _05432_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__a31o_1
X_14483_ clknet_leaf_6_clk _00997_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13503_ sha256cu.K\[27\] _06713_ _06718_ _00055_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__a22o_1
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ sha256cu.msg_scheduler.mreg_10\[24\] _04601_ VGND VGND VPWR VPWR _04605_
+ sky130_fd_sc_hd__or2_1
X_13434_ _03288_ _06722_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__and2_1
XFILLER_139_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10577_ sha256cu.msg_scheduler.mreg_8\[26\] _04554_ _04565_ _04557_ VGND VGND VPWR
+ VPWR _00742_ sky130_fd_sc_hd__o211a_1
XFILLER_10_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13365_ _06683_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_102_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_115_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12316_ _06101_ _06102_ _06105_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__o21a_1
XFILLER_54_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13296_ _06647_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ sha256cu.iter_processing.w\[27\] _05894_ _06052_ _05866_ VGND VGND VPWR VPWR
+ _00925_ sky130_fd_sc_hd__o211a_1
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12178_ sha256cu.data_in_padd\[24\] _05667_ _05986_ _05445_ VGND VGND VPWR VPWR _05987_
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11129_ _04769_ _04975_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__nor2_1
XFILLER_77_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14819_ clknet_leaf_104_clk _01333_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_08340_ _02943_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__or2_1
XFILLER_149_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08271_ _02332_ _02876_ _02877_ _02000_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__o211a_1
X_07222_ _01631_ _01879_ _01880_ _01883_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__a31o_1
XFILLER_118_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07153_ _01667_ _01640_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__nand2_1
XFILLER_145_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07084_ _01694_ _01762_ _01620_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07986_ _02599_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__inv_2
XFILLER_86_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09725_ _01973_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__buf_2
X_06937_ _01581_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__nor2_1
XFILLER_28_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09656_ sha256cu.m_out_digest.h_in\[20\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[20\]
+ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__a22o_1
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06868_ state\[3\] state\[2\] net257 VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__o21ba_1
X_08607_ sha256cu.m_out_digest.b_in\[25\] _03177_ _03176_ sha256cu.m_out_digest.a_in\[25\]
+ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__o22a_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06799_ net230 net233 net232 net236 VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__or4_2
X_09587_ sha256cu.m_out_digest.f_in\[27\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[27\]
+ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__o22a_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08538_ _03095_ _03113_ _03137_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__o21ba_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _03033_ _03034_ _03070_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__a21o_1
XFILLER_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10500_ sha256cu.msg_scheduler.mreg_7\[25\] _04513_ _04521_ _04516_ VGND VGND VPWR
+ VPWR _00709_ sky130_fd_sc_hd__o211a_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11480_ sha256cu.m_pad_pars.block_512\[36\]\[0\] _05304_ _05311_ _05322_ VGND VGND
+ VPWR VPWR _05323_ sky130_fd_sc_hd__a211o_1
XFILLER_136_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10431_ sha256cu.msg_scheduler.mreg_6\[27\] _04474_ _04482_ _04477_ VGND VGND VPWR
+ VPWR _00679_ sky130_fd_sc_hd__o211a_1
XFILLER_109_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10362_ sha256cu.msg_scheduler.mreg_6\[30\] _04441_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__or2_1
XFILLER_128_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13150_ _06569_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10293_ sha256cu.msg_scheduler.mreg_5\[0\] _04393_ _04403_ _04397_ VGND VGND VPWR
+ VPWR _00620_ sky130_fd_sc_hd__o211a_1
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12101_ _05911_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__or2_1
X_13081_ _06532_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12032_ sha256cu.msg_scheduler.mreg_9\[19\] sha256cu.msg_scheduler.mreg_0\[19\] VGND
+ VGND VPWR VPWR _05846_ sky130_fd_sc_hd__nand2_1
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13983_ clknet_leaf_55_clk _00529_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12934_ sha256cu.m_pad_pars.block_512\[34\]\[1\] _06453_ VGND VGND VPWR VPWR _06455_
+ sky130_fd_sc_hd__and2_1
XFILLER_19_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12865_ sha256cu.m_pad_pars.block_512\[30\]\[1\] _06416_ VGND VGND VPWR VPWR _06418_
+ sky130_fd_sc_hd__and2_1
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _01994_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__clkbuf_4
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ clknet_leaf_14_clk _01118_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12796_ _06381_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__clkbuf_1
X_11747_ sha256cu.msg_scheduler.mreg_1\[14\] sha256cu.msg_scheduler.mreg_1\[10\] VGND
+ VGND VPWR VPWR _05573_ sky130_fd_sc_hd__xnor2_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ clknet_leaf_8_clk _01049_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11678_ _05494_ _05496_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__nand2_1
X_14466_ clknet_leaf_101_clk _00980_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10629_ sha256cu.msg_scheduler.mreg_9\[16\] _04594_ _04595_ _04584_ VGND VGND VPWR
+ VPWR _00764_ sky130_fd_sc_hd__o211a_1
X_14397_ clknet_leaf_48_clk _00911_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[13\]
+ sky130_fd_sc_hd__dfxtp_4
X_13417_ sha256cu.m_pad_pars.block_512\[62\]\[5\] _01928_ VGND VGND VPWR VPWR _06710_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13348_ _06674_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__clkbuf_1
X_13279_ _06638_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07840_ _02455_ _02457_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07771_ _02349_ _02351_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__nor2_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09510_ _03951_ _03954_ _03981_ _02065_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__a31o_1
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09441_ _03914_ _03915_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09372_ _03846_ _03847_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__and2_1
X_08323_ sha256cu.m_out_digest.a_in\[27\] _02927_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08254_ sha256cu.iter_processing.w\[23\] _02860_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__xor2_1
XFILLER_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08185_ _02737_ _02755_ _02793_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__a21bo_1
X_07205_ _01804_ _01868_ _01644_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07136_ _01705_ _01808_ _01809_ _01598_ _01571_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__o221a_1
XFILLER_118_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07067_ _01649_ _01602_ _01694_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__or3_1
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07969_ _02583_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__inv_2
X_09708_ _04053_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__clkbuf_2
XFILLER_74_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10980_ sha256cu.m_pad_pars.block_512\[39\]\[1\] _04800_ _04826_ sha256cu.m_pad_pars.block_512\[51\]\[1\]
+ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__a22o_1
X_09639_ sha256cu.m_out_digest.h_in\[5\] _04037_ _04036_ sha256cu.m_out_digest.g_in\[5\]
+ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__a22o_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12650_ _06303_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__clkbuf_1
X_11601_ sha256cu.msg_scheduler.mreg_9\[0\] sha256cu.msg_scheduler.mreg_0\[0\] VGND
+ VGND VPWR VPWR _05434_ sky130_fd_sc_hd__nand2_1
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12581_ _06266_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14320_ clknet_leaf_90_clk _00014_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11532_ sha256cu.m_pad_pars.block_512\[16\]\[5\] _05285_ _05296_ sha256cu.m_pad_pars.block_512\[28\]\[5\]
+ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__a22o_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14251_ clknet_leaf_25_clk _00797_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11463_ _01935_ _05297_ _05305_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__and3_2
X_10414_ sha256cu.msg_scheduler.mreg_6\[20\] _04461_ _04472_ _04464_ VGND VGND VPWR
+ VPWR _00672_ sky130_fd_sc_hd__o211a_1
X_14182_ clknet_leaf_28_clk _00728_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ _06597_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13133_ _06560_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__clkbuf_1
X_11394_ _04768_ _05154_ _05237_ sha256cu.m_pad_pars.block_512\[5\]\[7\] VGND VGND
+ VPWR VPWR _05238_ sky130_fd_sc_hd__o22a_1
X_10345_ sha256cu.msg_scheduler.mreg_6\[23\] _04428_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__or2_1
XFILLER_151_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10276_ _04314_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__buf_2
XFILLER_3_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _06523_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__clkbuf_1
X_12015_ _05828_ _05829_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__and2_1
XFILLER_105_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13966_ clknet_leaf_55_clk _00512_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[20\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13897_ clknet_leaf_23_clk _00443_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12917_ sha256cu.m_pad_pars.block_512\[33\]\[1\] _06444_ VGND VGND VPWR VPWR _06446_
+ sky130_fd_sc_hd__and2_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12848_ sha256cu.m_pad_pars.block_512\[29\]\[1\] _06407_ VGND VGND VPWR VPWR _06409_
+ sky130_fd_sc_hd__and2_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12779_ _06372_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__clkbuf_1
X_14518_ clknet_leaf_114_clk _01032_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14449_ clknet_leaf_7_clk _00963_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09990_ sha256cu.msg_scheduler.mreg_0\[30\] _04221_ _04230_ _04224_ VGND VGND VPWR
+ VPWR _00490_ sky130_fd_sc_hd__o211a_1
XFILLER_115_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08941_ sha256cu.iter_processing.w\[10\] _02374_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__nand2_1
XFILLER_69_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08872_ _02332_ _03364_ _03365_ _03366_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__o211a_1
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07823_ _02332_ _02438_ _02441_ _02000_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__o211a_1
X_07754_ sha256cu.m_out_digest.g_in\[10\] sha256cu.m_out_digest.f_in\[10\] sha256cu.m_out_digest.e_in\[10\]
+ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__mux2_1
X_07685_ sha256cu.m_out_digest.h_in\[8\] _02306_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__xnor2_2
XFILLER_65_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09424_ sha256cu.m_out_digest.h_in\[27\] sha256cu.m_out_digest.d_in\[27\] VGND VGND
+ VPWR VPWR _03899_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_91_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09355_ _03830_ _03831_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__or2_1
XFILLER_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09286_ sha256cu.iter_processing.w\[22\] _02819_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__and2_1
X_08306_ _02909_ _02911_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08237_ _02069_ _02844_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__nor2_1
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08168_ sha256cu.m_out_digest.e_in\[27\] _02776_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__xnor2_4
XFILLER_4_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08099_ sha256cu.iter_processing.w\[19\] _02709_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__xnor2_1
X_07119_ _01631_ _01788_ _01789_ _01791_ _01794_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__a32o_1
X_10130_ sha256cu.msg_scheduler.mreg_2\[26\] _04301_ _04310_ _04304_ VGND VGND VPWR
+ VPWR _00550_ sky130_fd_sc_hd__o211a_1
XFILLER_122_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10061_ sha256cu.msg_scheduler.mreg_2\[29\] _04268_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__or2_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13820_ clknet_leaf_48_clk _00366_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_14\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_56_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13751_ clknet_leaf_63_clk _00297_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10963_ _04746_ _04758_ _04761_ _04807_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__o22a_1
XFILLER_16_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_43_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12702_ sha256cu.m_pad_pars.block_512\[20\]\[5\] _06325_ VGND VGND VPWR VPWR _06331_
+ sky130_fd_sc_hd__and2_1
X_13682_ clknet_leaf_66_clk _00228_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10894_ _04699_ _04760_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__nand2_2
X_12633_ _06294_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12564_ _06257_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__clkbuf_1
X_11515_ _05347_ _05349_ _05354_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__or3_2
X_14303_ clknet_leaf_95_clk _00027_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__dfxtp_1
X_14234_ clknet_leaf_19_clk _00780_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12495_ sha256cu.m_pad_pars.block_512\[8\]\[5\] _06214_ VGND VGND VPWR VPWR _06220_
+ sky130_fd_sc_hd__and2_1
X_11446_ sha256cu.m_pad_pars.block_512\[16\]\[0\] _05285_ _05288_ sha256cu.m_pad_pars.block_512\[48\]\[0\]
+ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__a22o_1
X_14165_ clknet_leaf_34_clk _00711_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11377_ sha256cu.m_pad_pars.block_512\[25\]\[6\] _05140_ _05141_ sha256cu.m_pad_pars.block_512\[29\]\[6\]
+ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__a22o_1
X_14096_ clknet_leaf_33_clk _00642_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10328_ _04396_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__buf_2
XFILLER_140_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13116_ _06551_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__clkbuf_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _06514_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__clkbuf_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ sha256cu.msg_scheduler.mreg_5\[18\] _04374_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__or2_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13949_ clknet_leaf_54_clk _00495_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[3\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_73_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07470_ _02032_ _02060_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__and2_1
XFILLER_22_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09140_ _03623_ _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__nor2_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09071_ sha256cu.m_out_digest.e_in\[14\] _02732_ _03557_ _03558_ _01913_ VGND VGND
+ VPWR VPWR _00237_ sky130_fd_sc_hd__a221o_1
X_08022_ _02594_ _02595_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__and2b_1
XFILLER_115_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09973_ sha256cu.msg_scheduler.mreg_0\[23\] _04208_ _04220_ _04211_ VGND VGND VPWR
+ VPWR _00483_ sky130_fd_sc_hd__o211a_1
XFILLER_104_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08924_ _03388_ _03391_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__o21a_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08855_ sha256cu.m_out_digest.h_in\[7\] sha256cu.m_out_digest.d_in\[7\] VGND VGND
+ VPWR VPWR _03350_ sky130_fd_sc_hd__nand2_1
XFILLER_111_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07806_ _02422_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__xnor2_2
X_08786_ _03240_ _03254_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__a21boi_2
XFILLER_85_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07737_ _02314_ _02312_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_64_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_53_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07668_ _02249_ _02251_ _02256_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__o21ai_1
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07599_ sha256cu.m_out_digest.b_in\[6\] sha256cu.m_out_digest.a_in\[6\] sha256cu.m_out_digest.c_in\[6\]
+ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a21o_1
XFILLER_111_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09407_ _03848_ _03856_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09338_ _02895_ _03815_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__xor2_1
XFILLER_40_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09269_ _03711_ _03728_ _03748_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__a21o_1
X_11300_ _04824_ _05004_ _05136_ _01952_ _05150_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__o221a_2
XFILLER_107_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12280_ _06058_ _06061_ _06057_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__a21boi_1
XFILLER_134_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11231_ _05081_ _04960_ _05082_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__o21a_1
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11162_ sha256cu.m_pad_pars.block_512\[2\]\[1\] _04999_ _04996_ sha256cu.m_pad_pars.block_512\[34\]\[1\]
+ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__a22o_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10113_ sha256cu.msg_scheduler.mreg_2\[19\] _04288_ _04300_ _04291_ VGND VGND VPWR
+ VPWR _00543_ sky130_fd_sc_hd__o211a_1
XFILLER_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11093_ _04725_ _04721_ _04951_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__or3b_1
XFILLER_0_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10044_ sha256cu.msg_scheduler.mreg_2\[22\] _04254_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__or2_1
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14921_ clknet_leaf_11_clk _01435_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14852_ clknet_leaf_100_clk _01366_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13803_ clknet_leaf_70_clk _00349_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_55_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
X_11995_ _05783_ _05788_ _05810_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__and3_1
XFILLER_91_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14783_ clknet_leaf_106_clk _01297_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[45\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13734_ clknet_leaf_81_clk _00280_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10946_ sha256cu.m_pad_pars.block_512\[11\]\[0\] _04790_ _04800_ sha256cu.m_pad_pars.block_512\[39\]\[0\]
+ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a221o_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13665_ clknet_leaf_85_clk _00211_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10877_ _04743_ sha256cu.m_pad_pars.add_512_block\[4\] VGND VGND VPWR VPWR _04744_
+ sky130_fd_sc_hd__nand2_2
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12616_ _06285_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13596_ clknet_leaf_68_clk _00142_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12547_ _06247_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _01479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12478_ sha256cu.m_pad_pars.block_512\[7\]\[5\] _06205_ VGND VGND VPWR VPWR _06211_
+ sky130_fd_sc_hd__and2_1
X_14217_ clknet_leaf_28_clk _00763_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11429_ _01985_ _05134_ _05266_ _05272_ _01970_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__a311o_1
XFILLER_153_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14148_ clknet_leaf_33_clk _00694_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ clknet_leaf_36_clk _00625_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ _01601_ _01589_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__or2_2
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08640_ sha256cu.m_out_digest.c_in\[20\] _03184_ _03182_ sha256cu.m_out_digest.b_in\[20\]
+ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__a22o_1
XFILLER_27_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
X_08571_ _03162_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__xnor2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07522_ _02104_ _02148_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07453_ sha256cu.m_out_digest.e_in\[27\] _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__xnor2_2
XFILLER_23_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09123_ _03553_ _03581_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__nand2_1
X_07384_ sha256cu.iter_processing.temp_case _01984_ _02006_ _02007_ VGND VGND VPWR
+ VPWR _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09054_ sha256cu.iter_processing.w\[14\] _02521_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__and2_1
XFILLER_135_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08005_ _02589_ _02590_ _02618_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__a21oi_2
XFILLER_116_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09956_ sha256cu.msg_scheduler.mreg_0\[15\] _04208_ _04210_ _04211_ VGND VGND VPWR
+ VPWR _00475_ sky130_fd_sc_hd__o211a_1
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08907_ _02302_ _03369_ _03370_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__a21boi_1
XFILLER_112_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09887_ sha256cu.msg_scheduler.mreg_12\[27\] _04167_ _04169_ _04157_ VGND VGND VPWR
+ VPWR _00442_ sky130_fd_sc_hd__o211a_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _03303_ _03301_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__or2b_1
XFILLER_18_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_122_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08769_ _03265_ _03266_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__nand2_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_404 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _05603_ _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__or2_1
X_10800_ _01566_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__buf_4
X_10731_ _04547_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__clkbuf_2
XFILLER_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13450_ _06730_ _06733_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__and2_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10662_ _04547_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__clkbuf_2
X_12401_ _06170_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10593_ sha256cu.msg_scheduler.mreg_10\[1\] _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__or2_1
X_13381_ _06691_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12332_ sha256cu.m_pad_pars.add_512_block\[1\] _01939_ _01947_ VGND VGND VPWR VPWR
+ _06132_ sky130_fd_sc_hd__and3_1
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12263_ _06066_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__nand2_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14002_ clknet_leaf_40_clk _00548_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11214_ sha256cu.m_pad_pars.block_512\[34\]\[5\] _04996_ _04981_ sha256cu.m_pad_pars.block_512\[54\]\[5\]
+ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__a22o_1
XFILLER_5_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12194_ _06000_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__nand2_1
XFILLER_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11145_ _04704_ _04993_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__or2_2
X_11076_ sha256cu.m_pad_pars.block_512\[39\]\[7\] _04795_ _04797_ VGND VGND VPWR VPWR
+ _04936_ sky130_fd_sc_hd__o21a_1
Xinput140 hash[225] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
X_10027_ sha256cu.msg_scheduler.mreg_1\[14\] _04247_ _04251_ _04250_ VGND VGND VPWR
+ VPWR _00506_ sky130_fd_sc_hd__o211a_1
Xinput151 hash[235] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput162 hash[245] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
X_14904_ clknet_leaf_125_clk _01418_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput184 hash[34] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_2
Xinput173 hash[255] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput195 hash[44] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_28_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_64_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14835_ clknet_leaf_0_clk _01349_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11978_ _05775_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__nand2_1
X_14766_ clknet_leaf_113_clk _01280_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13717_ clknet_leaf_65_clk _00263_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10929_ _04703_ _04771_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__or2_1
X_14697_ clknet_leaf_7_clk _01211_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13648_ clknet_leaf_51_clk _00194_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13579_ clknet_leaf_78_clk _00125_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09810_ sha256cu.msg_scheduler.mreg_14\[27\] _04120_ VGND VGND VPWR VPWR _04125_
+ sky130_fd_sc_hd__or2_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09741_ sha256cu.msg_scheduler.mreg_14\[29\] _04073_ _04085_ _04077_ VGND VGND VPWR
+ VPWR _00380_ sky130_fd_sc_hd__o211a_1
X_06953_ _01573_ _01642_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__nand2_2
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09672_ _01566_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__clkbuf_4
X_06884_ _01573_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__nand2_4
X_08623_ sha256cu.m_out_digest.c_in\[7\] _03179_ _03178_ sha256cu.m_out_digest.b_in\[7\]
+ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_19_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08554_ sha256cu.m_out_digest.h_in\[30\] _03116_ _03152_ VGND VGND VPWR VPWR _03153_
+ sky130_fd_sc_hd__a21oi_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _02127_ _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__xnor2_1
X_08485_ _03083_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__xor2_1
XFILLER_23_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07436_ _01911_ _02064_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__nor2_8
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07367_ sha256cu.m_pad_pars.add_out0\[6\] _01963_ _01998_ _02002_ VGND VGND VPWR
+ VPWR _02003_ sky130_fd_sc_hd__a31o_1
XFILLER_10_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09106_ _03590_ _03591_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__or2_1
XFILLER_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09037_ _03489_ _03505_ _03524_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__a21o_1
X_07298_ _01940_ _01941_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__nor2_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09939_ sha256cu.msg_scheduler.mreg_0\[8\] _04195_ _04201_ _04198_ VGND VGND VPWR
+ VPWR _00468_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12950_ _06463_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__clkbuf_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ sha256cu.msg_scheduler.mreg_14\[23\] sha256cu.msg_scheduler.mreg_14\[0\]
+ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12881_ _06426_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_201 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_212 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _05651_ _05653_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__or2_1
XFILLER_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_234 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14620_ clknet_leaf_122_clk _01134_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[24\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_245 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_267 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14551_ clknet_leaf_119_clk _01065_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11763_ _05585_ _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__xnor2_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10714_ sha256cu.msg_scheduler.mreg_10\[21\] _04633_ _04643_ _04636_ VGND VGND VPWR
+ VPWR _00801_ sky130_fd_sc_hd__o211a_1
X_11694_ _05521_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__nand2_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ clknet_leaf_6_clk _00996_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13502_ _06765_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_1
X_10645_ sha256cu.msg_scheduler.mreg_9\[23\] _04594_ _04604_ _04597_ VGND VGND VPWR
+ VPWR _00771_ sky130_fd_sc_hd__o211a_1
X_13433_ sha256cu.K\[1\] _06714_ _06719_ _00047_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__a22o_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13364_ sha256cu.m_pad_pars.block_512\[59\]\[3\] _06682_ VGND VGND VPWR VPWR _06683_
+ sky130_fd_sc_hd__and2_1
XFILLER_127_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10576_ sha256cu.msg_scheduler.mreg_9\[26\] _04561_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__or2_1
X_12315_ sha256cu.iter_processing.w\[30\] _05894_ _06117_ _01974_ VGND VGND VPWR VPWR
+ _00928_ sky130_fd_sc_hd__o211a_1
XFILLER_142_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13295_ sha256cu.m_pad_pars.block_512\[55\]\[2\] _06644_ VGND VGND VPWR VPWR _06647_
+ sky130_fd_sc_hd__and2_1
XFILLER_114_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12246_ _05442_ _06049_ _06050_ _06051_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__a31o_1
X_12177_ _05967_ _05984_ _05985_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__o21a_1
XFILLER_123_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11128_ _04725_ _04721_ _04720_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__or3_2
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11059_ _04779_ _04917_ _04918_ sha256cu.m_pad_pars.block_512\[47\]\[7\] VGND VGND
+ VPWR VPWR _04919_ sky130_fd_sc_hd__o22a_1
XFILLER_37_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14818_ clknet_leaf_104_clk _01332_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[49\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14749_ clknet_leaf_122_clk _01263_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[40\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08270_ sha256cu.m_out_digest.a_in\[23\] _02440_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__or2_1
XFILLER_20_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07221_ _00456_ _01881_ _01882_ _01663_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__o211a_1
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07152_ _01652_ _01819_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__nor2_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
X_07083_ _01643_ _01602_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__nand2_1
XFILLER_114_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07985_ sha256cu.m_out_digest.e_in\[27\] _02598_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__xnor2_2
XFILLER_75_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09724_ sha256cu.iter_processing.w\[22\] _04067_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__or2_1
X_06936_ _01588_ _01626_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__or2_1
X_09655_ sha256cu.m_out_digest.h_in\[19\] _04041_ _04040_ sha256cu.m_out_digest.g_in\[19\]
+ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__a22o_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06867_ _01562_ _01563_ net257 VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08606_ sha256cu.m_out_digest.b_in\[24\] _03177_ _03176_ _02083_ VGND VGND VPWR VPWR
+ _00151_ sky130_fd_sc_hd__o22a_1
XFILLER_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09586_ sha256cu.m_out_digest.f_in\[26\] _04029_ _04028_ sha256cu.m_out_digest.e_in\[26\]
+ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__a22o_1
X_06798_ _01492_ _01493_ _01494_ _01495_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__or4_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08537_ _03134_ _03136_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ _03068_ _03069_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__nand2_1
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07419_ _02046_ _02047_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__and2b_1
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10430_ sha256cu.msg_scheduler.mreg_7\[27\] _04481_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__or2_1
XFILLER_109_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08399_ _02999_ _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10361_ sha256cu.msg_scheduler.mreg_5\[29\] _04434_ _04442_ _04437_ VGND VGND VPWR
+ VPWR _00649_ sky130_fd_sc_hd__o211a_1
XFILLER_128_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10292_ sha256cu.msg_scheduler.mreg_6\[0\] _04401_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__or2_1
X_12100_ _05883_ _05891_ _05910_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__and3_1
X_13080_ sha256cu.m_pad_pars.block_512\[42\]\[6\] _06525_ VGND VGND VPWR VPWR _06532_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12031_ sha256cu.msg_scheduler.mreg_9\[19\] sha256cu.msg_scheduler.mreg_0\[19\] VGND
+ VGND VPWR VPWR _05845_ sky130_fd_sc_hd__or2_1
XFILLER_151_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13982_ clknet_leaf_55_clk _00528_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12933_ _06454_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _06417_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ sha256cu.data_in_padd\[9\] _05448_ _05638_ _05463_ VGND VGND VPWR VPWR _05639_
+ sky130_fd_sc_hd__a211o_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ clknet_leaf_14_clk _01117_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[22\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12795_ sha256cu.m_pad_pars.block_512\[26\]\[0\] _06380_ VGND VGND VPWR VPWR _06381_
+ sky130_fd_sc_hd__and2_1
X_11746_ _05570_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__nand2_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14534_ clknet_leaf_102_clk _01048_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _05497_ _05499_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__or2_1
X_14465_ clknet_leaf_99_clk _00979_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10628_ sha256cu.msg_scheduler.mreg_10\[16\] _04588_ VGND VGND VPWR VPWR _04595_
+ sky130_fd_sc_hd__or2_1
X_14396_ clknet_leaf_47_clk _00910_ VGND VGND VPWR VPWR sha256cu.iter_processing.w\[12\]
+ sky130_fd_sc_hd__dfxtp_4
X_13416_ _06709_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10559_ sha256cu.msg_scheduler.mreg_8\[18\] _04554_ _04555_ _04543_ VGND VGND VPWR
+ VPWR _00734_ sky130_fd_sc_hd__o211a_1
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13347_ sha256cu.m_pad_pars.block_512\[58\]\[3\] _06671_ VGND VGND VPWR VPWR _06674_
+ sky130_fd_sc_hd__and2_1
X_13278_ sha256cu.m_pad_pars.block_512\[54\]\[2\] _06635_ VGND VGND VPWR VPWR _06638_
+ sky130_fd_sc_hd__and2_1
X_12229_ _06033_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nand2_1
XFILLER_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07770_ _02378_ _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__xor2_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09440_ _03877_ _03881_ _03875_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__o21a_1
XFILLER_52_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09371_ _03846_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__nor2_1
XFILLER_18_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08322_ _02084_ sha256cu.m_out_digest.a_in\[6\] VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08253_ _02858_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07204_ _01593_ _01646_ _01750_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__and3_1
XFILLER_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08184_ _02754_ _02752_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__or2b_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07135_ _01578_ _01612_ _01640_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07066_ _01590_ _01733_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__nand2_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07968_ _02555_ _02556_ _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__nand3_2
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09707_ sha256cu.msg_scheduler.mreg_14\[14\] _04060_ _04066_ _04064_ VGND VGND VPWR
+ VPWR _00365_ sky130_fd_sc_hd__o211a_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_06919_ _01592_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07899_ _02481_ _02479_ _02513_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__o31a_1
XFILLER_83_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09638_ sha256cu.m_out_digest.h_in\[4\] _04039_ _04038_ sha256cu.m_out_digest.g_in\[4\]
+ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__o22a_1
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09569_ sha256cu.m_out_digest.f_in\[11\] _04027_ _04026_ sha256cu.m_out_digest.e_in\[11\]
+ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__o22a_1
XFILLER_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11600_ _05432_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__clkbuf_4
X_12580_ sha256cu.m_pad_pars.block_512\[13\]\[4\] _06261_ VGND VGND VPWR VPWR _06266_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11531_ sha256cu.m_pad_pars.block_512\[44\]\[5\] _05298_ _05320_ sha256cu.m_pad_pars.block_512\[40\]\[5\]
+ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__a221o_1
XFILLER_128_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14250_ clknet_leaf_25_clk _00796_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_10\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11462_ _04792_ _05136_ _04909_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__o21a_1
X_10413_ sha256cu.msg_scheduler.mreg_7\[20\] _04468_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__or2_1
X_14181_ clknet_leaf_28_clk _00727_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_8\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11393_ _04954_ _01956_ _04786_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__and3b_1
X_13201_ sha256cu.m_pad_pars.block_512\[49\]\[6\] _06590_ VGND VGND VPWR VPWR _06597_
+ sky130_fd_sc_hd__and2_1
X_10344_ sha256cu.msg_scheduler.mreg_5\[22\] _04421_ _04432_ _04424_ VGND VGND VPWR
+ VPWR _00642_ sky130_fd_sc_hd__o211a_1
XFILLER_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13132_ sha256cu.m_pad_pars.block_512\[45\]\[6\] _06553_ VGND VGND VPWR VPWR _06560_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10275_ sha256cu.msg_scheduler.mreg_4\[25\] _04380_ _04392_ _04383_ VGND VGND VPWR
+ VPWR _00613_ sky130_fd_sc_hd__o211a_1
XFILLER_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ sha256cu.m_pad_pars.block_512\[41\]\[6\] _06516_ VGND VGND VPWR VPWR _06523_
+ sky130_fd_sc_hd__and2_1
X_12014_ _05826_ _05827_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__nand2_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13965_ clknet_leaf_57_clk _00511_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[19\]
+ sky130_fd_sc_hd__dfxtp_2
X_13896_ clknet_leaf_22_clk _00442_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12916_ _06445_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__clkbuf_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _06408_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12778_ sha256cu.m_pad_pars.block_512\[25\]\[0\] _06371_ VGND VGND VPWR VPWR _06372_
+ sky130_fd_sc_hd__and2_1
X_11729_ _05530_ _05534_ _05531_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__a21boi_1
X_14517_ clknet_leaf_3_clk _01031_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14448_ clknet_leaf_9_clk _00962_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_14379_ clknet_leaf_110_clk _00893_ VGND VGND VPWR VPWR sha256cu.data_in_padd\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08940_ sha256cu.iter_processing.w\[10\] _02374_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__or2_1
XFILLER_115_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08871_ _01973_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__clkbuf_8
XFILLER_111_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07822_ sha256cu.m_out_digest.a_in\[11\] _02440_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__or2_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07753_ sha256cu.m_out_digest.b_in\[10\] sha256cu.m_out_digest.a_in\[10\] sha256cu.m_out_digest.c_in\[10\]
+ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__a21o_1
X_07684_ _02304_ _02305_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__xnor2_4
X_09423_ _03885_ _03886_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__nand2_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09354_ _03830_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__nand2_1
X_08305_ sha256cu.iter_processing.w\[23\] _02860_ _02910_ VGND VGND VPWR VPWR _02911_
+ sky130_fd_sc_hd__a21oi_1
X_09285_ sha256cu.iter_processing.w\[22\] _02819_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__nor2_1
X_08236_ _02839_ _02843_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08167_ sha256cu.m_out_digest.e_in\[14\] sha256cu.m_out_digest.e_in\[0\] VGND VGND
+ VPWR VPWR _02776_ sky130_fd_sc_hd__xnor2_4
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07118_ _00456_ _01793_ _01629_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08098_ _02707_ _02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07049_ _01725_ _01731_ _01571_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__mux2_1
X_10060_ sha256cu.msg_scheduler.mreg_1\[28\] _04260_ _04270_ _04264_ VGND VGND VPWR
+ VPWR _00520_ sky130_fd_sc_hd__o211a_1
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13750_ clknet_leaf_65_clk _00296_ VGND VGND VPWR VPWR sha256cu.m_out_digest.g_in\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10962_ _01919_ _04736_ _04755_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__and3_2
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12701_ _06330_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13681_ clknet_leaf_66_clk _00227_ VGND VGND VPWR VPWR sha256cu.m_out_digest.e_in\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_44_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10893_ _04748_ _01940_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__nor2_2
X_12632_ sha256cu.m_pad_pars.block_512\[16\]\[4\] _06289_ VGND VGND VPWR VPWR _06294_
+ sky130_fd_sc_hd__and2_1
XFILLER_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12563_ sha256cu.m_pad_pars.block_512\[12\]\[4\] _06252_ VGND VGND VPWR VPWR _06257_
+ sky130_fd_sc_hd__and2_1
XFILLER_145_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12494_ _06219_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_1
X_14302_ clknet_4_5_0_clk _00026_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11514_ sha256cu.m_pad_pars.block_512\[0\]\[3\] _05314_ _05350_ _05353_ VGND VGND
+ VPWR VPWR _05354_ sky130_fd_sc_hd__a211o_1
X_14233_ clknet_leaf_19_clk _00779_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11445_ _04705_ _05286_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__o21a_2
XFILLER_152_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14164_ clknet_leaf_34_clk _00710_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11376_ sha256cu.m_pad_pars.block_512\[13\]\[6\] _05128_ _05144_ sha256cu.m_pad_pars.block_512\[9\]\[6\]
+ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__a22o_1
X_10327_ sha256cu.msg_scheduler.mreg_6\[15\] _04415_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__or2_1
X_14095_ clknet_leaf_33_clk _00641_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13115_ sha256cu.m_pad_pars.block_512\[44\]\[6\] _06544_ VGND VGND VPWR VPWR _06551_
+ sky130_fd_sc_hd__and2_1
X_10258_ sha256cu.msg_scheduler.mreg_4\[17\] _04380_ _04382_ _04383_ VGND VGND VPWR
+ VPWR _00605_ sky130_fd_sc_hd__o211a_1
XFILLER_140_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ sha256cu.m_pad_pars.block_512\[40\]\[6\] _06507_ VGND VGND VPWR VPWR _06514_
+ sky130_fd_sc_hd__and2_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10189_ sha256cu.msg_scheduler.mreg_3\[19\] _04341_ _04343_ _04344_ VGND VGND VPWR
+ VPWR _00575_ sky130_fd_sc_hd__o211a_1
XFILLER_79_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13948_ clknet_leaf_53_clk _00494_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_1\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13879_ clknet_leaf_20_clk _00425_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_12\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09070_ _03553_ _03556_ _02515_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__o21a_1
XFILLER_30_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08021_ _02592_ _02611_ _02633_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09972_ sha256cu.msg_scheduler.mreg_1\[23\] _04215_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__or2_1
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08923_ _03356_ _03367_ _03386_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__a21o_1
XFILLER_130_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08854_ sha256cu.m_out_digest.h_in\[7\] sha256cu.m_out_digest.d_in\[7\] VGND VGND
+ VPWR VPWR _03349_ sky130_fd_sc_hd__or2_1
X_07805_ _02381_ _02385_ _02423_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__o21a_1
X_08785_ _03253_ _03251_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__or2b_1
X_07736_ _02335_ _02356_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07667_ _02260_ _02289_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__xnor2_2
XFILLER_53_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07598_ sha256cu.m_out_digest.b_in\[6\] sha256cu.m_out_digest.a_in\[6\] VGND VGND
+ VPWR VPWR _02222_ sky130_fd_sc_hd__or2_1
XFILLER_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09406_ _03877_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__xor2_1
XFILLER_41_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09337_ _03813_ _03814_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__nand2_1
XFILLER_139_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09268_ _03711_ _03728_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__and3_1
X_08219_ _02824_ _02826_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__nor2_1
X_09199_ _03676_ _03680_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__and2_1
XFILLER_153_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11230_ _04698_ _04908_ _04785_ sha256cu.m_pad_pars.block_512\[26\]\[7\] VGND VGND
+ VPWR VPWR _05082_ sky130_fd_sc_hd__a31o_1
XFILLER_136_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11161_ sha256cu.m_pad_pars.block_512\[6\]\[1\] _04957_ _04964_ sha256cu.m_pad_pars.block_512\[26\]\[1\]
+ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__a22o_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10112_ sha256cu.msg_scheduler.mreg_3\[19\] _04295_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__or2_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11092_ sha256cu.m_pad_pars.add_out2\[3\] sha256cu.m_pad_pars.add_out2\[2\] VGND
+ VGND VPWR VPWR _04951_ sky130_fd_sc_hd__and2b_1
X_10043_ _04166_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__buf_2
XFILLER_75_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14920_ clknet_leaf_10_clk _01434_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[62\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14851_ clknet_leaf_98_clk _01365_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[53\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13802_ clknet_leaf_82_clk _00348_ VGND VGND VPWR VPWR sha256cu.m_out_digest.h_in\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11994_ _05807_ _05809_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14782_ clknet_leaf_123_clk _01296_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[44\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13733_ clknet_leaf_83_clk _00279_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10945_ sha256cu.m_pad_pars.block_512\[43\]\[0\] _04804_ _04811_ sha256cu.m_pad_pars.block_512\[31\]\[0\]
+ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__a22o_1
XFILLER_71_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13664_ clknet_leaf_84_clk _00210_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10876_ sha256cu.m_pad_pars.add_512_block\[5\] VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__inv_2
XFILLER_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12615_ sha256cu.m_pad_pars.block_512\[15\]\[4\] _06280_ VGND VGND VPWR VPWR _06285_
+ sky130_fd_sc_hd__and2_1
X_13595_ clknet_leaf_67_clk _00141_ VGND VGND VPWR VPWR sha256cu.m_out_digest.b_in\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12546_ sha256cu.m_pad_pars.block_512\[11\]\[5\] _06241_ VGND VGND VPWR VPWR _06247_
+ sky130_fd_sc_hd__and2_1
XFILLER_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12477_ _06210_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__clkbuf_1
X_14216_ clknet_leaf_28_clk _00762_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_9\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_4 _01479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11428_ _05125_ _05134_ _05267_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__a31o_1
XFILLER_153_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14147_ clknet_leaf_35_clk _00693_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_7\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11359_ sha256cu.m_pad_pars.block_512\[37\]\[4\] _05165_ _05205_ _05024_ VGND VGND
+ VPWR VPWR _05206_ sky130_fd_sc_hd__a22o_1
XFILLER_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14078_ clknet_leaf_36_clk _00624_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_5\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ sha256cu.m_pad_pars.block_512\[39\]\[6\] _06498_ VGND VGND VPWR VPWR _06505_
+ sky130_fd_sc_hd__and2_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08570_ _03163_ _03168_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07521_ _02145_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nand2_1
XFILLER_81_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07452_ sha256cu.m_out_digest.e_in\[13\] sha256cu.m_out_digest.e_in\[8\] VGND VGND
+ VPWR VPWR _02080_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07383_ _02014_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09122_ _03606_ _03607_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__and2_1
XFILLER_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09053_ sha256cu.iter_processing.w\[14\] _02521_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__nor2_1
XFILLER_151_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08004_ _02616_ _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__nand2_1
XFILLER_116_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09955_ _04116_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__clkbuf_4
XFILLER_106_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08906_ _02344_ _03398_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__xor2_1
XFILLER_100_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09886_ sha256cu.msg_scheduler.mreg_13\[27\] _04160_ VGND VGND VPWR VPWR _04169_
+ sky130_fd_sc_hd__or2_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _03331_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__xor2_1
XFILLER_106_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ sha256cu.m_out_digest.h_in\[4\] sha256cu.m_out_digest.d_in\[4\] VGND VGND
+ VPWR VPWR _03266_ sky130_fd_sc_hd__nand2_1
XANTENNA_405 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _02336_ _02337_ _02338_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__a21o_1
XFILLER_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08699_ _02024_ _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__xor2_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10730_ sha256cu.msg_scheduler.mreg_10\[28\] _04646_ _04652_ _04649_ VGND VGND VPWR
+ VPWR _00808_ sky130_fd_sc_hd__o211a_1
XFILLER_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10661_ sha256cu.msg_scheduler.mreg_9\[30\] _04607_ _04613_ _04610_ VGND VGND VPWR
+ VPWR _00778_ sky130_fd_sc_hd__o211a_1
X_12400_ sha256cu.m_pad_pars.block_512\[3\]\[0\] _06169_ VGND VGND VPWR VPWR _06170_
+ sky130_fd_sc_hd__and2_1
XFILLER_41_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10592_ _04547_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__clkbuf_2
X_13380_ sha256cu.m_pad_pars.block_512\[60\]\[3\] _06682_ VGND VGND VPWR VPWR _06691_
+ sky130_fd_sc_hd__and2_1
X_12331_ _06131_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12262_ sha256cu.msg_scheduler.mreg_14\[15\] sha256cu.msg_scheduler.mreg_14\[13\]
+ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__xor2_1
X_14001_ clknet_leaf_55_clk _00547_ VGND VGND VPWR VPWR sha256cu.msg_scheduler.mreg_2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11213_ sha256cu.m_pad_pars.block_512\[30\]\[5\] _05009_ _04977_ sha256cu.m_pad_pars.block_512\[46\]\[5\]
+ _05066_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__a221o_1
XFILLER_134_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12193_ _05998_ _05999_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or2_1
XFILLER_122_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11144_ sha256cu.m_pad_pars.block_512\[14\]\[0\] _04989_ _04996_ sha256cu.m_pad_pars.block_512\[34\]\[0\]
+ _05002_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a221o_1
XFILLER_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11075_ _04758_ _04933_ _04934_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__o21ba_1
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput163 hash[246] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xinput141 hash[226] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlymetal6s2s_1
X_10026_ sha256cu.msg_scheduler.mreg_2\[14\] _04241_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__or2_1
Xinput152 hash[236] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xinput130 hash[216] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14903_ clknet_leaf_124_clk _01417_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[60\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput196 hash[45] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput185 hash[35] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
Xinput174 hash[25] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_4
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14834_ clknet_leaf_2_clk _01348_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[51\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11977_ _05792_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__and2_1
X_14765_ clknet_leaf_16_clk _01279_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[42\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13716_ clknet_leaf_61_clk _00262_ VGND VGND VPWR VPWR sha256cu.m_out_digest.f_in\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10928_ _04770_ _04794_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__nor2_2
XFILLER_149_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14696_ clknet_leaf_7_clk _01210_ VGND VGND VPWR VPWR sha256cu.m_pad_pars.block_512\[34\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13647_ clknet_leaf_73_clk _00193_ VGND VGND VPWR VPWR sha256cu.m_out_digest.d_in\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10859_ _01979_ _04730_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__nor2_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ clknet_leaf_78_clk _00124_ VGND VGND VPWR VPWR sha256cu.m_out_digest.a_in\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12529_ sha256cu.m_pad_pars.block_512\[10\]\[5\] _06232_ VGND VGND VPWR VPWR _06238_
+ sky130_fd_sc_hd__and2_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09740_ sha256cu.iter_processing.w\[29\] _04080_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__or2_1
X_06952_ _01577_ _01580_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__nand2_2
.ends

